module MulAddRecFNToRaw_postMul_1( // @[:chipyard.TestHarness.RocketConfig.fir@236971.2]
  input          io_fromPreMul_isSigNaNAny, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input          io_fromPreMul_isNaNAOrB, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input          io_fromPreMul_isInfA, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input          io_fromPreMul_isZeroA, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input          io_fromPreMul_isInfB, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input          io_fromPreMul_isZeroB, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input          io_fromPreMul_signProd, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input          io_fromPreMul_isNaNC, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input          io_fromPreMul_isInfC, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input          io_fromPreMul_isZeroC, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input  [12:0]  io_fromPreMul_sExpSum, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input          io_fromPreMul_doSubMags, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input          io_fromPreMul_CIsDominant, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input  [5:0]   io_fromPreMul_CDom_CAlignDist, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input  [54:0]  io_fromPreMul_highAlignedSigC, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input          io_fromPreMul_bit0AlignedSigC, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input  [106:0] io_mulAddResult, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  input  [2:0]   io_roundingMode, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  output         io_invalidExc, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  output         io_rawOut_isNaN, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  output         io_rawOut_isInf, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  output         io_rawOut_isZero, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  output         io_rawOut_sign, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  output [12:0]  io_rawOut_sExp, // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
  output [55:0]  io_rawOut_sig // @[:chipyard.TestHarness.RocketConfig.fir@236972.4]
);
  wire  roundingMode_min; // @[MulAddRecFN.scala 188:45:chipyard.TestHarness.RocketConfig.fir@236975.4]
  wire  CDom_sign; // @[MulAddRecFN.scala 192:42:chipyard.TestHarness.RocketConfig.fir@236976.4]
  wire [54:0] _T_2; // @[MulAddRecFN.scala 195:47:chipyard.TestHarness.RocketConfig.fir@236979.4]
  wire [54:0] _T_3; // @[MulAddRecFN.scala 194:16:chipyard.TestHarness.RocketConfig.fir@236980.4]
  wire [161:0] sigSum; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236983.4]
  wire [1:0] _T_6; // @[MulAddRecFN.scala 205:69:chipyard.TestHarness.RocketConfig.fir@236984.4]
  wire [12:0] _GEN_0; // @[MulAddRecFN.scala 205:43:chipyard.TestHarness.RocketConfig.fir@236985.4]
  wire [12:0] CDom_sExp; // @[MulAddRecFN.scala 205:43:chipyard.TestHarness.RocketConfig.fir@236987.4]
  wire [107:0] _T_10; // @[MulAddRecFN.scala 208:13:chipyard.TestHarness.RocketConfig.fir@236989.4]
  wire [107:0] _T_14; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236993.4]
  wire [107:0] CDom_absSigSum; // @[MulAddRecFN.scala 207:12:chipyard.TestHarness.RocketConfig.fir@236994.4]
  wire [52:0] _T_16; // @[MulAddRecFN.scala 217:14:chipyard.TestHarness.RocketConfig.fir@236996.4]
  wire  _T_17; // @[MulAddRecFN.scala 217:36:chipyard.TestHarness.RocketConfig.fir@236997.4]
  wire  _T_19; // @[MulAddRecFN.scala 218:37:chipyard.TestHarness.RocketConfig.fir@236999.4]
  wire  CDom_absSigSumExtra; // @[MulAddRecFN.scala 216:12:chipyard.TestHarness.RocketConfig.fir@237000.4]
  wire [170:0] _GEN_1; // @[MulAddRecFN.scala 221:24:chipyard.TestHarness.RocketConfig.fir@237001.4]
  wire [170:0] _T_20; // @[MulAddRecFN.scala 221:24:chipyard.TestHarness.RocketConfig.fir@237001.4]
  wire [57:0] CDom_mainSig; // @[MulAddRecFN.scala 221:56:chipyard.TestHarness.RocketConfig.fir@237002.4]
  wire [54:0] _T_22; // @[MulAddRecFN.scala 224:53:chipyard.TestHarness.RocketConfig.fir@237004.4]
  wire  _T_25; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237008.4]
  wire  _T_27; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237011.4]
  wire  _T_29; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237014.4]
  wire  _T_31; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237017.4]
  wire  _T_33; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237020.4]
  wire  _T_35; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237023.4]
  wire  _T_37; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237026.4]
  wire  _T_39; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237029.4]
  wire  _T_41; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237032.4]
  wire  _T_43; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237035.4]
  wire  _T_45; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237038.4]
  wire  _T_47; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237041.4]
  wire  _T_49; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237044.4]
  wire  _T_51; // @[primitives.scala 124:57:chipyard.TestHarness.RocketConfig.fir@237047.4]
  wire [6:0] _T_57; // @[primitives.scala 125:20:chipyard.TestHarness.RocketConfig.fir@237054.4]
  wire [13:0] _T_64; // @[primitives.scala 125:20:chipyard.TestHarness.RocketConfig.fir@237061.4]
  wire [3:0] _T_66; // @[primitives.scala 51:21:chipyard.TestHarness.RocketConfig.fir@237063.4]
  wire [16:0] _T_67; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@237064.4]
  wire [7:0] _T_73; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237070.4]
  wire [7:0] _T_75; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237072.4]
  wire [7:0] _T_77; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237074.4]
  wire [7:0] _T_78; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237075.4]
  wire [7:0] _GEN_2; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237080.4]
  wire [7:0] _T_83; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237080.4]
  wire [7:0] _T_85; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237082.4]
  wire [7:0] _T_87; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237084.4]
  wire [7:0] _T_88; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237085.4]
  wire [7:0] _GEN_3; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237090.4]
  wire [7:0] _T_93; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237090.4]
  wire [7:0] _T_95; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237092.4]
  wire [7:0] _T_97; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237094.4]
  wire [7:0] _T_98; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237095.4]
  wire [12:0] _T_112; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237109.4]
  wire [13:0] _GEN_4; // @[MulAddRecFN.scala 224:72:chipyard.TestHarness.RocketConfig.fir@237110.4]
  wire [13:0] _T_113; // @[MulAddRecFN.scala 224:72:chipyard.TestHarness.RocketConfig.fir@237110.4]
  wire  CDom_reduced4SigExtra; // @[MulAddRecFN.scala 225:73:chipyard.TestHarness.RocketConfig.fir@237111.4]
  wire  _T_116; // @[MulAddRecFN.scala 228:32:chipyard.TestHarness.RocketConfig.fir@237114.4]
  wire  _T_117; // @[MulAddRecFN.scala 228:36:chipyard.TestHarness.RocketConfig.fir@237115.4]
  wire  _T_118; // @[MulAddRecFN.scala 228:61:chipyard.TestHarness.RocketConfig.fir@237116.4]
  wire [55:0] CDom_sig; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237117.4]
  wire  notCDom_signSigSum; // @[MulAddRecFN.scala 234:36:chipyard.TestHarness.RocketConfig.fir@237118.4]
  wire [108:0] _T_120; // @[MulAddRecFN.scala 237:13:chipyard.TestHarness.RocketConfig.fir@237120.4]
  wire [108:0] _GEN_5; // @[MulAddRecFN.scala 238:41:chipyard.TestHarness.RocketConfig.fir@237122.4]
  wire [108:0] _T_123; // @[MulAddRecFN.scala 238:41:chipyard.TestHarness.RocketConfig.fir@237123.4]
  wire [108:0] notCDom_absSigSum; // @[MulAddRecFN.scala 236:12:chipyard.TestHarness.RocketConfig.fir@237124.4]
  wire  _T_126; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237128.4]
  wire  _T_128; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237131.4]
  wire  _T_130; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237134.4]
  wire  _T_132; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237137.4]
  wire  _T_134; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237140.4]
  wire  _T_136; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237143.4]
  wire  _T_138; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237146.4]
  wire  _T_140; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237149.4]
  wire  _T_142; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237152.4]
  wire  _T_144; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237155.4]
  wire  _T_146; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237158.4]
  wire  _T_148; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237161.4]
  wire  _T_150; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237164.4]
  wire  _T_152; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237167.4]
  wire  _T_154; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237170.4]
  wire  _T_156; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237173.4]
  wire  _T_158; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237176.4]
  wire  _T_160; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237179.4]
  wire  _T_162; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237182.4]
  wire  _T_164; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237185.4]
  wire  _T_166; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237188.4]
  wire  _T_168; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237191.4]
  wire  _T_170; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237194.4]
  wire  _T_172; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237197.4]
  wire  _T_174; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237200.4]
  wire  _T_176; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237203.4]
  wire  _T_178; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237206.4]
  wire  _T_180; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237209.4]
  wire  _T_182; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237212.4]
  wire  _T_184; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237215.4]
  wire  _T_186; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237218.4]
  wire  _T_188; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237221.4]
  wire  _T_190; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237224.4]
  wire  _T_192; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237227.4]
  wire  _T_194; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237230.4]
  wire  _T_196; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237233.4]
  wire  _T_198; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237236.4]
  wire  _T_200; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237239.4]
  wire  _T_202; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237242.4]
  wire  _T_204; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237245.4]
  wire  _T_206; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237248.4]
  wire  _T_208; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237251.4]
  wire  _T_210; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237254.4]
  wire  _T_212; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237257.4]
  wire  _T_214; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237260.4]
  wire  _T_216; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237263.4]
  wire  _T_218; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237266.4]
  wire  _T_220; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237269.4]
  wire  _T_222; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237272.4]
  wire  _T_224; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237275.4]
  wire  _T_226; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237278.4]
  wire  _T_228; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237281.4]
  wire  _T_230; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237284.4]
  wire  _T_232; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237287.4]
  wire  _T_234; // @[primitives.scala 107:57:chipyard.TestHarness.RocketConfig.fir@237290.4]
  wire [5:0] _T_239; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237296.4]
  wire [12:0] _T_246; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237303.4]
  wire [6:0] _T_252; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237309.4]
  wire [26:0] _T_260; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237317.4]
  wire [6:0] _T_266; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237323.4]
  wire [13:0] _T_273; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237330.4]
  wire [6:0] _T_279; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237336.4]
  wire [54:0] notCDom_reduced2AbsSigSum; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237345.4]
  wire [5:0] _T_343; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237401.4]
  wire [5:0] _T_344; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237402.4]
  wire [5:0] _T_345; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237403.4]
  wire [5:0] _T_346; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237404.4]
  wire [5:0] _T_347; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237405.4]
  wire [5:0] _T_348; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237406.4]
  wire [5:0] _T_349; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237407.4]
  wire [5:0] _T_350; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237408.4]
  wire [5:0] _T_351; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237409.4]
  wire [5:0] _T_352; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237410.4]
  wire [5:0] _T_353; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237411.4]
  wire [5:0] _T_354; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237412.4]
  wire [5:0] _T_355; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237413.4]
  wire [5:0] _T_356; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237414.4]
  wire [5:0] _T_357; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237415.4]
  wire [5:0] _T_358; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237416.4]
  wire [5:0] _T_359; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237417.4]
  wire [5:0] _T_360; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237418.4]
  wire [5:0] _T_361; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237419.4]
  wire [5:0] _T_362; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237420.4]
  wire [5:0] _T_363; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237421.4]
  wire [5:0] _T_364; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237422.4]
  wire [5:0] _T_365; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237423.4]
  wire [5:0] _T_366; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237424.4]
  wire [5:0] _T_367; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237425.4]
  wire [5:0] _T_368; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237426.4]
  wire [5:0] _T_369; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237427.4]
  wire [5:0] _T_370; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237428.4]
  wire [5:0] _T_371; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237429.4]
  wire [5:0] _T_372; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237430.4]
  wire [5:0] _T_373; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237431.4]
  wire [5:0] _T_374; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237432.4]
  wire [5:0] _T_375; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237433.4]
  wire [5:0] _T_376; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237434.4]
  wire [5:0] _T_377; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237435.4]
  wire [5:0] _T_378; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237436.4]
  wire [5:0] _T_379; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237437.4]
  wire [5:0] _T_380; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237438.4]
  wire [5:0] _T_381; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237439.4]
  wire [5:0] _T_382; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237440.4]
  wire [5:0] _T_383; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237441.4]
  wire [5:0] _T_384; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237442.4]
  wire [5:0] _T_385; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237443.4]
  wire [5:0] _T_386; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237444.4]
  wire [5:0] _T_387; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237445.4]
  wire [5:0] _T_388; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237446.4]
  wire [5:0] _T_389; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237447.4]
  wire [5:0] _T_390; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237448.4]
  wire [5:0] _T_391; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237449.4]
  wire [5:0] _T_392; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237450.4]
  wire [5:0] _T_393; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237451.4]
  wire [5:0] _T_394; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237452.4]
  wire [5:0] _T_395; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237453.4]
  wire [5:0] notCDom_normDistReduced2; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237454.4]
  wire [6:0] notCDom_nearNormDist; // @[MulAddRecFN.scala 242:56:chipyard.TestHarness.RocketConfig.fir@237455.4]
  wire [7:0] _T_396; // @[MulAddRecFN.scala 243:69:chipyard.TestHarness.RocketConfig.fir@237456.4]
  wire [12:0] _GEN_6; // @[MulAddRecFN.scala 243:46:chipyard.TestHarness.RocketConfig.fir@237457.4]
  wire [12:0] notCDom_sExp; // @[MulAddRecFN.scala 243:46:chipyard.TestHarness.RocketConfig.fir@237459.4]
  wire [235:0] _GEN_7; // @[MulAddRecFN.scala 245:27:chipyard.TestHarness.RocketConfig.fir@237460.4]
  wire [235:0] _T_399; // @[MulAddRecFN.scala 245:27:chipyard.TestHarness.RocketConfig.fir@237460.4]
  wire [57:0] notCDom_mainSig; // @[MulAddRecFN.scala 245:50:chipyard.TestHarness.RocketConfig.fir@237461.4]
  wire  _T_404; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237467.4]
  wire  _T_406; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237470.4]
  wire  _T_408; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237473.4]
  wire  _T_410; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237476.4]
  wire  _T_412; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237479.4]
  wire  _T_414; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237482.4]
  wire  _T_416; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237485.4]
  wire  _T_418; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237488.4]
  wire  _T_420; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237491.4]
  wire  _T_422; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237494.4]
  wire  _T_424; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237497.4]
  wire  _T_426; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237500.4]
  wire  _T_428; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237503.4]
  wire  _T_430; // @[primitives.scala 107:57:chipyard.TestHarness.RocketConfig.fir@237506.4]
  wire [6:0] _T_436; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237513.4]
  wire [13:0] _T_443; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237520.4]
  wire [4:0] _T_445; // @[primitives.scala 51:21:chipyard.TestHarness.RocketConfig.fir@237522.4]
  wire [32:0] _T_446; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@237523.4]
  wire [7:0] _T_452; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237529.4]
  wire [7:0] _T_454; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237531.4]
  wire [7:0] _T_456; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237533.4]
  wire [7:0] _T_457; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237534.4]
  wire [7:0] _GEN_8; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237539.4]
  wire [7:0] _T_462; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237539.4]
  wire [7:0] _T_464; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237541.4]
  wire [7:0] _T_466; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237543.4]
  wire [7:0] _T_467; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237544.4]
  wire [7:0] _GEN_9; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237549.4]
  wire [7:0] _T_472; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237549.4]
  wire [7:0] _T_474; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237551.4]
  wire [7:0] _T_476; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237553.4]
  wire [7:0] _T_477; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237554.4]
  wire [12:0] _T_491; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237568.4]
  wire [13:0] _GEN_10; // @[MulAddRecFN.scala 249:78:chipyard.TestHarness.RocketConfig.fir@237569.4]
  wire [13:0] _T_492; // @[MulAddRecFN.scala 249:78:chipyard.TestHarness.RocketConfig.fir@237569.4]
  wire  notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 251:11:chipyard.TestHarness.RocketConfig.fir@237570.4]
  wire  _T_495; // @[MulAddRecFN.scala 254:35:chipyard.TestHarness.RocketConfig.fir@237573.4]
  wire  _T_496; // @[MulAddRecFN.scala 254:39:chipyard.TestHarness.RocketConfig.fir@237574.4]
  wire [55:0] notCDom_sig; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237575.4]
  wire  notCDom_completeCancellation; // @[MulAddRecFN.scala 257:50:chipyard.TestHarness.RocketConfig.fir@237577.4]
  wire  _T_498; // @[MulAddRecFN.scala 261:36:chipyard.TestHarness.RocketConfig.fir@237578.4]
  wire  notCDom_sign; // @[MulAddRecFN.scala 259:12:chipyard.TestHarness.RocketConfig.fir@237579.4]
  wire  notNaN_isInfProd; // @[MulAddRecFN.scala 266:49:chipyard.TestHarness.RocketConfig.fir@237580.4]
  wire  notNaN_isInfOut; // @[MulAddRecFN.scala 267:44:chipyard.TestHarness.RocketConfig.fir@237581.4]
  wire  _T_499; // @[MulAddRecFN.scala 269:32:chipyard.TestHarness.RocketConfig.fir@237582.4]
  wire  notNaN_addZeros; // @[MulAddRecFN.scala 269:58:chipyard.TestHarness.RocketConfig.fir@237583.4]
  wire  _T_500; // @[MulAddRecFN.scala 274:31:chipyard.TestHarness.RocketConfig.fir@237584.4]
  wire  _T_501; // @[MulAddRecFN.scala 273:35:chipyard.TestHarness.RocketConfig.fir@237585.4]
  wire  _T_502; // @[MulAddRecFN.scala 275:32:chipyard.TestHarness.RocketConfig.fir@237586.4]
  wire  _T_503; // @[MulAddRecFN.scala 274:57:chipyard.TestHarness.RocketConfig.fir@237587.4]
  wire  _T_504; // @[MulAddRecFN.scala 276:10:chipyard.TestHarness.RocketConfig.fir@237588.4]
  wire  _T_506; // @[MulAddRecFN.scala 276:36:chipyard.TestHarness.RocketConfig.fir@237590.4]
  wire  _T_507; // @[MulAddRecFN.scala 277:61:chipyard.TestHarness.RocketConfig.fir@237591.4]
  wire  _T_508; // @[MulAddRecFN.scala 278:35:chipyard.TestHarness.RocketConfig.fir@237592.4]
  wire  _T_511; // @[MulAddRecFN.scala 285:14:chipyard.TestHarness.RocketConfig.fir@237598.4]
  wire  _T_512; // @[MulAddRecFN.scala 285:42:chipyard.TestHarness.RocketConfig.fir@237599.4]
  wire  _T_514; // @[MulAddRecFN.scala 287:27:chipyard.TestHarness.RocketConfig.fir@237602.4]
  wire  _T_515; // @[MulAddRecFN.scala 288:31:chipyard.TestHarness.RocketConfig.fir@237603.4]
  wire  _T_516; // @[MulAddRecFN.scala 287:54:chipyard.TestHarness.RocketConfig.fir@237604.4]
  wire  _T_517; // @[MulAddRecFN.scala 289:29:chipyard.TestHarness.RocketConfig.fir@237605.4]
  wire  _T_518; // @[MulAddRecFN.scala 289:26:chipyard.TestHarness.RocketConfig.fir@237606.4]
  wire  _T_519; // @[MulAddRecFN.scala 289:48:chipyard.TestHarness.RocketConfig.fir@237607.4]
  wire  _T_520; // @[MulAddRecFN.scala 290:36:chipyard.TestHarness.RocketConfig.fir@237608.4]
  wire  _T_521; // @[MulAddRecFN.scala 288:43:chipyard.TestHarness.RocketConfig.fir@237609.4]
  wire  _T_522; // @[MulAddRecFN.scala 291:26:chipyard.TestHarness.RocketConfig.fir@237610.4]
  wire  _T_523; // @[MulAddRecFN.scala 292:37:chipyard.TestHarness.RocketConfig.fir@237611.4]
  wire  _T_524; // @[MulAddRecFN.scala 291:46:chipyard.TestHarness.RocketConfig.fir@237612.4]
  wire  _T_525; // @[MulAddRecFN.scala 290:48:chipyard.TestHarness.RocketConfig.fir@237613.4]
  wire  _T_526; // @[MulAddRecFN.scala 293:10:chipyard.TestHarness.RocketConfig.fir@237614.4]
  wire  _T_527; // @[MulAddRecFN.scala 293:31:chipyard.TestHarness.RocketConfig.fir@237615.4]
  wire  _T_528; // @[MulAddRecFN.scala 293:28:chipyard.TestHarness.RocketConfig.fir@237616.4]
  wire  _T_529; // @[MulAddRecFN.scala 294:17:chipyard.TestHarness.RocketConfig.fir@237617.4]
  wire  _T_530; // @[MulAddRecFN.scala 293:49:chipyard.TestHarness.RocketConfig.fir@237618.4]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[MulAddRecFN.scala 188:45:chipyard.TestHarness.RocketConfig.fir@236975.4]
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42:chipyard.TestHarness.RocketConfig.fir@236976.4]
  assign _T_2 = io_fromPreMul_highAlignedSigC + 55'h1; // @[MulAddRecFN.scala 195:47:chipyard.TestHarness.RocketConfig.fir@236979.4]
  assign _T_3 = io_mulAddResult[106] ? _T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16:chipyard.TestHarness.RocketConfig.fir@236980.4]
  assign sigSum = {_T_3,io_mulAddResult[105:0],io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236983.4]
  assign _T_6 = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69:chipyard.TestHarness.RocketConfig.fir@236984.4]
  assign _GEN_0 = {{11{_T_6[1]}},_T_6}; // @[MulAddRecFN.scala 205:43:chipyard.TestHarness.RocketConfig.fir@236985.4]
  assign CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43:chipyard.TestHarness.RocketConfig.fir@236987.4]
  assign _T_10 = ~sigSum[161:54]; // @[MulAddRecFN.scala 208:13:chipyard.TestHarness.RocketConfig.fir@236989.4]
  assign _T_14 = {1'h0,io_fromPreMul_highAlignedSigC[54:53],sigSum[159:55]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236993.4]
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? _T_10 : _T_14; // @[MulAddRecFN.scala 207:12:chipyard.TestHarness.RocketConfig.fir@236994.4]
  assign _T_16 = ~sigSum[53:1]; // @[MulAddRecFN.scala 217:14:chipyard.TestHarness.RocketConfig.fir@236996.4]
  assign _T_17 = |_T_16; // @[MulAddRecFN.scala 217:36:chipyard.TestHarness.RocketConfig.fir@236997.4]
  assign _T_19 = |sigSum[54:1]; // @[MulAddRecFN.scala 218:37:chipyard.TestHarness.RocketConfig.fir@236999.4]
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _T_17 : _T_19; // @[MulAddRecFN.scala 216:12:chipyard.TestHarness.RocketConfig.fir@237000.4]
  assign _GEN_1 = {{63'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24:chipyard.TestHarness.RocketConfig.fir@237001.4]
  assign _T_20 = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24:chipyard.TestHarness.RocketConfig.fir@237001.4]
  assign CDom_mainSig = _T_20[107:50]; // @[MulAddRecFN.scala 221:56:chipyard.TestHarness.RocketConfig.fir@237002.4]
  assign _T_22 = {CDom_absSigSum[52:0], 2'h0}; // @[MulAddRecFN.scala 224:53:chipyard.TestHarness.RocketConfig.fir@237004.4]
  assign _T_25 = |_T_22[3:0]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237008.4]
  assign _T_27 = |_T_22[7:4]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237011.4]
  assign _T_29 = |_T_22[11:8]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237014.4]
  assign _T_31 = |_T_22[15:12]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237017.4]
  assign _T_33 = |_T_22[19:16]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237020.4]
  assign _T_35 = |_T_22[23:20]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237023.4]
  assign _T_37 = |_T_22[27:24]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237026.4]
  assign _T_39 = |_T_22[31:28]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237029.4]
  assign _T_41 = |_T_22[35:32]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237032.4]
  assign _T_43 = |_T_22[39:36]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237035.4]
  assign _T_45 = |_T_22[43:40]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237038.4]
  assign _T_47 = |_T_22[47:44]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237041.4]
  assign _T_49 = |_T_22[51:48]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@237044.4]
  assign _T_51 = |_T_22[54:52]; // @[primitives.scala 124:57:chipyard.TestHarness.RocketConfig.fir@237047.4]
  assign _T_57 = {_T_37,_T_35,_T_33,_T_31,_T_29,_T_27,_T_25}; // @[primitives.scala 125:20:chipyard.TestHarness.RocketConfig.fir@237054.4]
  assign _T_64 = {_T_51,_T_49,_T_47,_T_45,_T_43,_T_41,_T_39,_T_57}; // @[primitives.scala 125:20:chipyard.TestHarness.RocketConfig.fir@237061.4]
  assign _T_66 = ~io_fromPreMul_CDom_CAlignDist[5:2]; // @[primitives.scala 51:21:chipyard.TestHarness.RocketConfig.fir@237063.4]
  assign _T_67 = -17'sh10000 >>> _T_66; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@237064.4]
  assign _T_73 = {{4'd0}, _T_67[8:5]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237070.4]
  assign _T_75 = {_T_67[4:1], 4'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237072.4]
  assign _T_77 = _T_75 & 8'hf0; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237074.4]
  assign _T_78 = _T_73 | _T_77; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237075.4]
  assign _GEN_2 = {{2'd0}, _T_78[7:2]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237080.4]
  assign _T_83 = _GEN_2 & 8'h33; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237080.4]
  assign _T_85 = {_T_78[5:0], 2'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237082.4]
  assign _T_87 = _T_85 & 8'hcc; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237084.4]
  assign _T_88 = _T_83 | _T_87; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237085.4]
  assign _GEN_3 = {{1'd0}, _T_88[7:1]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237090.4]
  assign _T_93 = _GEN_3 & 8'h55; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237090.4]
  assign _T_95 = {_T_88[6:0], 1'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237092.4]
  assign _T_97 = _T_95 & 8'haa; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237094.4]
  assign _T_98 = _T_93 | _T_97; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237095.4]
  assign _T_112 = {_T_98,_T_67[9],_T_67[10],_T_67[11],_T_67[12],_T_67[13]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237109.4]
  assign _GEN_4 = {{1'd0}, _T_112}; // @[MulAddRecFN.scala 224:72:chipyard.TestHarness.RocketConfig.fir@237110.4]
  assign _T_113 = _T_64 & _GEN_4; // @[MulAddRecFN.scala 224:72:chipyard.TestHarness.RocketConfig.fir@237110.4]
  assign CDom_reduced4SigExtra = |_T_113; // @[MulAddRecFN.scala 225:73:chipyard.TestHarness.RocketConfig.fir@237111.4]
  assign _T_116 = |CDom_mainSig[2:0]; // @[MulAddRecFN.scala 228:32:chipyard.TestHarness.RocketConfig.fir@237114.4]
  assign _T_117 = _T_116 | CDom_reduced4SigExtra; // @[MulAddRecFN.scala 228:36:chipyard.TestHarness.RocketConfig.fir@237115.4]
  assign _T_118 = _T_117 | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61:chipyard.TestHarness.RocketConfig.fir@237116.4]
  assign CDom_sig = {CDom_mainSig[57:3],_T_118}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237117.4]
  assign notCDom_signSigSum = sigSum[109]; // @[MulAddRecFN.scala 234:36:chipyard.TestHarness.RocketConfig.fir@237118.4]
  assign _T_120 = ~sigSum[108:0]; // @[MulAddRecFN.scala 237:13:chipyard.TestHarness.RocketConfig.fir@237120.4]
  assign _GEN_5 = {{108'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41:chipyard.TestHarness.RocketConfig.fir@237122.4]
  assign _T_123 = sigSum[108:0] + _GEN_5; // @[MulAddRecFN.scala 238:41:chipyard.TestHarness.RocketConfig.fir@237123.4]
  assign notCDom_absSigSum = notCDom_signSigSum ? _T_120 : _T_123; // @[MulAddRecFN.scala 236:12:chipyard.TestHarness.RocketConfig.fir@237124.4]
  assign _T_126 = |notCDom_absSigSum[1:0]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237128.4]
  assign _T_128 = |notCDom_absSigSum[3:2]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237131.4]
  assign _T_130 = |notCDom_absSigSum[5:4]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237134.4]
  assign _T_132 = |notCDom_absSigSum[7:6]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237137.4]
  assign _T_134 = |notCDom_absSigSum[9:8]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237140.4]
  assign _T_136 = |notCDom_absSigSum[11:10]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237143.4]
  assign _T_138 = |notCDom_absSigSum[13:12]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237146.4]
  assign _T_140 = |notCDom_absSigSum[15:14]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237149.4]
  assign _T_142 = |notCDom_absSigSum[17:16]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237152.4]
  assign _T_144 = |notCDom_absSigSum[19:18]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237155.4]
  assign _T_146 = |notCDom_absSigSum[21:20]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237158.4]
  assign _T_148 = |notCDom_absSigSum[23:22]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237161.4]
  assign _T_150 = |notCDom_absSigSum[25:24]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237164.4]
  assign _T_152 = |notCDom_absSigSum[27:26]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237167.4]
  assign _T_154 = |notCDom_absSigSum[29:28]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237170.4]
  assign _T_156 = |notCDom_absSigSum[31:30]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237173.4]
  assign _T_158 = |notCDom_absSigSum[33:32]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237176.4]
  assign _T_160 = |notCDom_absSigSum[35:34]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237179.4]
  assign _T_162 = |notCDom_absSigSum[37:36]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237182.4]
  assign _T_164 = |notCDom_absSigSum[39:38]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237185.4]
  assign _T_166 = |notCDom_absSigSum[41:40]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237188.4]
  assign _T_168 = |notCDom_absSigSum[43:42]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237191.4]
  assign _T_170 = |notCDom_absSigSum[45:44]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237194.4]
  assign _T_172 = |notCDom_absSigSum[47:46]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237197.4]
  assign _T_174 = |notCDom_absSigSum[49:48]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237200.4]
  assign _T_176 = |notCDom_absSigSum[51:50]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237203.4]
  assign _T_178 = |notCDom_absSigSum[53:52]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237206.4]
  assign _T_180 = |notCDom_absSigSum[55:54]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237209.4]
  assign _T_182 = |notCDom_absSigSum[57:56]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237212.4]
  assign _T_184 = |notCDom_absSigSum[59:58]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237215.4]
  assign _T_186 = |notCDom_absSigSum[61:60]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237218.4]
  assign _T_188 = |notCDom_absSigSum[63:62]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237221.4]
  assign _T_190 = |notCDom_absSigSum[65:64]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237224.4]
  assign _T_192 = |notCDom_absSigSum[67:66]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237227.4]
  assign _T_194 = |notCDom_absSigSum[69:68]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237230.4]
  assign _T_196 = |notCDom_absSigSum[71:70]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237233.4]
  assign _T_198 = |notCDom_absSigSum[73:72]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237236.4]
  assign _T_200 = |notCDom_absSigSum[75:74]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237239.4]
  assign _T_202 = |notCDom_absSigSum[77:76]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237242.4]
  assign _T_204 = |notCDom_absSigSum[79:78]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237245.4]
  assign _T_206 = |notCDom_absSigSum[81:80]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237248.4]
  assign _T_208 = |notCDom_absSigSum[83:82]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237251.4]
  assign _T_210 = |notCDom_absSigSum[85:84]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237254.4]
  assign _T_212 = |notCDom_absSigSum[87:86]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237257.4]
  assign _T_214 = |notCDom_absSigSum[89:88]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237260.4]
  assign _T_216 = |notCDom_absSigSum[91:90]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237263.4]
  assign _T_218 = |notCDom_absSigSum[93:92]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237266.4]
  assign _T_220 = |notCDom_absSigSum[95:94]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237269.4]
  assign _T_222 = |notCDom_absSigSum[97:96]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237272.4]
  assign _T_224 = |notCDom_absSigSum[99:98]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237275.4]
  assign _T_226 = |notCDom_absSigSum[101:100]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237278.4]
  assign _T_228 = |notCDom_absSigSum[103:102]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237281.4]
  assign _T_230 = |notCDom_absSigSum[105:104]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237284.4]
  assign _T_232 = |notCDom_absSigSum[107:106]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237287.4]
  assign _T_234 = |notCDom_absSigSum[108]; // @[primitives.scala 107:57:chipyard.TestHarness.RocketConfig.fir@237290.4]
  assign _T_239 = {_T_136,_T_134,_T_132,_T_130,_T_128,_T_126}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237296.4]
  assign _T_246 = {_T_150,_T_148,_T_146,_T_144,_T_142,_T_140,_T_138,_T_239}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237303.4]
  assign _T_252 = {_T_164,_T_162,_T_160,_T_158,_T_156,_T_154,_T_152}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237309.4]
  assign _T_260 = {_T_178,_T_176,_T_174,_T_172,_T_170,_T_168,_T_166,_T_252,_T_246}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237317.4]
  assign _T_266 = {_T_192,_T_190,_T_188,_T_186,_T_184,_T_182,_T_180}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237323.4]
  assign _T_273 = {_T_206,_T_204,_T_202,_T_200,_T_198,_T_196,_T_194,_T_266}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237330.4]
  assign _T_279 = {_T_220,_T_218,_T_216,_T_214,_T_212,_T_210,_T_208}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237336.4]
  assign notCDom_reduced2AbsSigSum = {_T_234,_T_232,_T_230,_T_228,_T_226,_T_224,_T_222,_T_279,_T_273,_T_260}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237345.4]
  assign _T_343 = notCDom_reduced2AbsSigSum[1] ? 6'h35 : 6'h36; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237401.4]
  assign _T_344 = notCDom_reduced2AbsSigSum[2] ? 6'h34 : _T_343; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237402.4]
  assign _T_345 = notCDom_reduced2AbsSigSum[3] ? 6'h33 : _T_344; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237403.4]
  assign _T_346 = notCDom_reduced2AbsSigSum[4] ? 6'h32 : _T_345; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237404.4]
  assign _T_347 = notCDom_reduced2AbsSigSum[5] ? 6'h31 : _T_346; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237405.4]
  assign _T_348 = notCDom_reduced2AbsSigSum[6] ? 6'h30 : _T_347; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237406.4]
  assign _T_349 = notCDom_reduced2AbsSigSum[7] ? 6'h2f : _T_348; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237407.4]
  assign _T_350 = notCDom_reduced2AbsSigSum[8] ? 6'h2e : _T_349; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237408.4]
  assign _T_351 = notCDom_reduced2AbsSigSum[9] ? 6'h2d : _T_350; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237409.4]
  assign _T_352 = notCDom_reduced2AbsSigSum[10] ? 6'h2c : _T_351; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237410.4]
  assign _T_353 = notCDom_reduced2AbsSigSum[11] ? 6'h2b : _T_352; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237411.4]
  assign _T_354 = notCDom_reduced2AbsSigSum[12] ? 6'h2a : _T_353; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237412.4]
  assign _T_355 = notCDom_reduced2AbsSigSum[13] ? 6'h29 : _T_354; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237413.4]
  assign _T_356 = notCDom_reduced2AbsSigSum[14] ? 6'h28 : _T_355; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237414.4]
  assign _T_357 = notCDom_reduced2AbsSigSum[15] ? 6'h27 : _T_356; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237415.4]
  assign _T_358 = notCDom_reduced2AbsSigSum[16] ? 6'h26 : _T_357; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237416.4]
  assign _T_359 = notCDom_reduced2AbsSigSum[17] ? 6'h25 : _T_358; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237417.4]
  assign _T_360 = notCDom_reduced2AbsSigSum[18] ? 6'h24 : _T_359; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237418.4]
  assign _T_361 = notCDom_reduced2AbsSigSum[19] ? 6'h23 : _T_360; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237419.4]
  assign _T_362 = notCDom_reduced2AbsSigSum[20] ? 6'h22 : _T_361; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237420.4]
  assign _T_363 = notCDom_reduced2AbsSigSum[21] ? 6'h21 : _T_362; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237421.4]
  assign _T_364 = notCDom_reduced2AbsSigSum[22] ? 6'h20 : _T_363; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237422.4]
  assign _T_365 = notCDom_reduced2AbsSigSum[23] ? 6'h1f : _T_364; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237423.4]
  assign _T_366 = notCDom_reduced2AbsSigSum[24] ? 6'h1e : _T_365; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237424.4]
  assign _T_367 = notCDom_reduced2AbsSigSum[25] ? 6'h1d : _T_366; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237425.4]
  assign _T_368 = notCDom_reduced2AbsSigSum[26] ? 6'h1c : _T_367; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237426.4]
  assign _T_369 = notCDom_reduced2AbsSigSum[27] ? 6'h1b : _T_368; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237427.4]
  assign _T_370 = notCDom_reduced2AbsSigSum[28] ? 6'h1a : _T_369; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237428.4]
  assign _T_371 = notCDom_reduced2AbsSigSum[29] ? 6'h19 : _T_370; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237429.4]
  assign _T_372 = notCDom_reduced2AbsSigSum[30] ? 6'h18 : _T_371; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237430.4]
  assign _T_373 = notCDom_reduced2AbsSigSum[31] ? 6'h17 : _T_372; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237431.4]
  assign _T_374 = notCDom_reduced2AbsSigSum[32] ? 6'h16 : _T_373; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237432.4]
  assign _T_375 = notCDom_reduced2AbsSigSum[33] ? 6'h15 : _T_374; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237433.4]
  assign _T_376 = notCDom_reduced2AbsSigSum[34] ? 6'h14 : _T_375; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237434.4]
  assign _T_377 = notCDom_reduced2AbsSigSum[35] ? 6'h13 : _T_376; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237435.4]
  assign _T_378 = notCDom_reduced2AbsSigSum[36] ? 6'h12 : _T_377; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237436.4]
  assign _T_379 = notCDom_reduced2AbsSigSum[37] ? 6'h11 : _T_378; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237437.4]
  assign _T_380 = notCDom_reduced2AbsSigSum[38] ? 6'h10 : _T_379; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237438.4]
  assign _T_381 = notCDom_reduced2AbsSigSum[39] ? 6'hf : _T_380; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237439.4]
  assign _T_382 = notCDom_reduced2AbsSigSum[40] ? 6'he : _T_381; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237440.4]
  assign _T_383 = notCDom_reduced2AbsSigSum[41] ? 6'hd : _T_382; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237441.4]
  assign _T_384 = notCDom_reduced2AbsSigSum[42] ? 6'hc : _T_383; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237442.4]
  assign _T_385 = notCDom_reduced2AbsSigSum[43] ? 6'hb : _T_384; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237443.4]
  assign _T_386 = notCDom_reduced2AbsSigSum[44] ? 6'ha : _T_385; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237444.4]
  assign _T_387 = notCDom_reduced2AbsSigSum[45] ? 6'h9 : _T_386; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237445.4]
  assign _T_388 = notCDom_reduced2AbsSigSum[46] ? 6'h8 : _T_387; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237446.4]
  assign _T_389 = notCDom_reduced2AbsSigSum[47] ? 6'h7 : _T_388; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237447.4]
  assign _T_390 = notCDom_reduced2AbsSigSum[48] ? 6'h6 : _T_389; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237448.4]
  assign _T_391 = notCDom_reduced2AbsSigSum[49] ? 6'h5 : _T_390; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237449.4]
  assign _T_392 = notCDom_reduced2AbsSigSum[50] ? 6'h4 : _T_391; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237450.4]
  assign _T_393 = notCDom_reduced2AbsSigSum[51] ? 6'h3 : _T_392; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237451.4]
  assign _T_394 = notCDom_reduced2AbsSigSum[52] ? 6'h2 : _T_393; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237452.4]
  assign _T_395 = notCDom_reduced2AbsSigSum[53] ? 6'h1 : _T_394; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237453.4]
  assign notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[54] ? 6'h0 : _T_395; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@237454.4]
  assign notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56:chipyard.TestHarness.RocketConfig.fir@237455.4]
  assign _T_396 = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69:chipyard.TestHarness.RocketConfig.fir@237456.4]
  assign _GEN_6 = {{5{_T_396[7]}},_T_396}; // @[MulAddRecFN.scala 243:46:chipyard.TestHarness.RocketConfig.fir@237457.4]
  assign notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_6); // @[MulAddRecFN.scala 243:46:chipyard.TestHarness.RocketConfig.fir@237459.4]
  assign _GEN_7 = {{127'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27:chipyard.TestHarness.RocketConfig.fir@237460.4]
  assign _T_399 = _GEN_7 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27:chipyard.TestHarness.RocketConfig.fir@237460.4]
  assign notCDom_mainSig = _T_399[109:52]; // @[MulAddRecFN.scala 245:50:chipyard.TestHarness.RocketConfig.fir@237461.4]
  assign _T_404 = |notCDom_reduced2AbsSigSum[1:0]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237467.4]
  assign _T_406 = |notCDom_reduced2AbsSigSum[3:2]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237470.4]
  assign _T_408 = |notCDom_reduced2AbsSigSum[5:4]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237473.4]
  assign _T_410 = |notCDom_reduced2AbsSigSum[7:6]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237476.4]
  assign _T_412 = |notCDom_reduced2AbsSigSum[9:8]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237479.4]
  assign _T_414 = |notCDom_reduced2AbsSigSum[11:10]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237482.4]
  assign _T_416 = |notCDom_reduced2AbsSigSum[13:12]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237485.4]
  assign _T_418 = |notCDom_reduced2AbsSigSum[15:14]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237488.4]
  assign _T_420 = |notCDom_reduced2AbsSigSum[17:16]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237491.4]
  assign _T_422 = |notCDom_reduced2AbsSigSum[19:18]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237494.4]
  assign _T_424 = |notCDom_reduced2AbsSigSum[21:20]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237497.4]
  assign _T_426 = |notCDom_reduced2AbsSigSum[23:22]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237500.4]
  assign _T_428 = |notCDom_reduced2AbsSigSum[25:24]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@237503.4]
  assign _T_430 = |notCDom_reduced2AbsSigSum[26]; // @[primitives.scala 107:57:chipyard.TestHarness.RocketConfig.fir@237506.4]
  assign _T_436 = {_T_416,_T_414,_T_412,_T_410,_T_408,_T_406,_T_404}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237513.4]
  assign _T_443 = {_T_430,_T_428,_T_426,_T_424,_T_422,_T_420,_T_418,_T_436}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@237520.4]
  assign _T_445 = ~notCDom_normDistReduced2[5:1]; // @[primitives.scala 51:21:chipyard.TestHarness.RocketConfig.fir@237522.4]
  assign _T_446 = -33'sh100000000 >>> _T_445; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@237523.4]
  assign _T_452 = {{4'd0}, _T_446[8:5]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237529.4]
  assign _T_454 = {_T_446[4:1], 4'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237531.4]
  assign _T_456 = _T_454 & 8'hf0; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237533.4]
  assign _T_457 = _T_452 | _T_456; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237534.4]
  assign _GEN_8 = {{2'd0}, _T_457[7:2]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237539.4]
  assign _T_462 = _GEN_8 & 8'h33; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237539.4]
  assign _T_464 = {_T_457[5:0], 2'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237541.4]
  assign _T_466 = _T_464 & 8'hcc; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237543.4]
  assign _T_467 = _T_462 | _T_466; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237544.4]
  assign _GEN_9 = {{1'd0}, _T_467[7:1]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237549.4]
  assign _T_472 = _GEN_9 & 8'h55; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237549.4]
  assign _T_474 = {_T_467[6:0], 1'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237551.4]
  assign _T_476 = _T_474 & 8'haa; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237553.4]
  assign _T_477 = _T_472 | _T_476; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237554.4]
  assign _T_491 = {_T_477,_T_446[9],_T_446[10],_T_446[11],_T_446[12],_T_446[13]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237568.4]
  assign _GEN_10 = {{1'd0}, _T_491}; // @[MulAddRecFN.scala 249:78:chipyard.TestHarness.RocketConfig.fir@237569.4]
  assign _T_492 = _T_443 & _GEN_10; // @[MulAddRecFN.scala 249:78:chipyard.TestHarness.RocketConfig.fir@237569.4]
  assign notCDom_reduced4SigExtra = |_T_492; // @[MulAddRecFN.scala 251:11:chipyard.TestHarness.RocketConfig.fir@237570.4]
  assign _T_495 = |notCDom_mainSig[2:0]; // @[MulAddRecFN.scala 254:35:chipyard.TestHarness.RocketConfig.fir@237573.4]
  assign _T_496 = _T_495 | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39:chipyard.TestHarness.RocketConfig.fir@237574.4]
  assign notCDom_sig = {notCDom_mainSig[57:3],_T_496}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237575.4]
  assign notCDom_completeCancellation = notCDom_sig[55:54] == 2'h0; // @[MulAddRecFN.scala 257:50:chipyard.TestHarness.RocketConfig.fir@237577.4]
  assign _T_498 = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36:chipyard.TestHarness.RocketConfig.fir@237578.4]
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : _T_498; // @[MulAddRecFN.scala 259:12:chipyard.TestHarness.RocketConfig.fir@237579.4]
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49:chipyard.TestHarness.RocketConfig.fir@237580.4]
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44:chipyard.TestHarness.RocketConfig.fir@237581.4]
  assign _T_499 = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 269:32:chipyard.TestHarness.RocketConfig.fir@237582.4]
  assign notNaN_addZeros = _T_499 & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58:chipyard.TestHarness.RocketConfig.fir@237583.4]
  assign _T_500 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31:chipyard.TestHarness.RocketConfig.fir@237584.4]
  assign _T_501 = io_fromPreMul_isSigNaNAny | _T_500; // @[MulAddRecFN.scala 273:35:chipyard.TestHarness.RocketConfig.fir@237585.4]
  assign _T_502 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32:chipyard.TestHarness.RocketConfig.fir@237586.4]
  assign _T_503 = _T_501 | _T_502; // @[MulAddRecFN.scala 274:57:chipyard.TestHarness.RocketConfig.fir@237587.4]
  assign _T_504 = ~io_fromPreMul_isNaNAOrB; // @[MulAddRecFN.scala 276:10:chipyard.TestHarness.RocketConfig.fir@237588.4]
  assign _T_506 = _T_504 & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36:chipyard.TestHarness.RocketConfig.fir@237590.4]
  assign _T_507 = _T_506 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61:chipyard.TestHarness.RocketConfig.fir@237591.4]
  assign _T_508 = _T_507 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35:chipyard.TestHarness.RocketConfig.fir@237592.4]
  assign _T_511 = ~io_fromPreMul_CIsDominant; // @[MulAddRecFN.scala 285:14:chipyard.TestHarness.RocketConfig.fir@237598.4]
  assign _T_512 = _T_511 & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42:chipyard.TestHarness.RocketConfig.fir@237599.4]
  assign _T_514 = notNaN_isInfProd & io_fromPreMul_signProd; // @[MulAddRecFN.scala 287:27:chipyard.TestHarness.RocketConfig.fir@237602.4]
  assign _T_515 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31:chipyard.TestHarness.RocketConfig.fir@237603.4]
  assign _T_516 = _T_514 | _T_515; // @[MulAddRecFN.scala 287:54:chipyard.TestHarness.RocketConfig.fir@237604.4]
  assign _T_517 = ~roundingMode_min; // @[MulAddRecFN.scala 289:29:chipyard.TestHarness.RocketConfig.fir@237605.4]
  assign _T_518 = notNaN_addZeros & _T_517; // @[MulAddRecFN.scala 289:26:chipyard.TestHarness.RocketConfig.fir@237606.4]
  assign _T_519 = _T_518 & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48:chipyard.TestHarness.RocketConfig.fir@237607.4]
  assign _T_520 = _T_519 & CDom_sign; // @[MulAddRecFN.scala 290:36:chipyard.TestHarness.RocketConfig.fir@237608.4]
  assign _T_521 = _T_516 | _T_520; // @[MulAddRecFN.scala 288:43:chipyard.TestHarness.RocketConfig.fir@237609.4]
  assign _T_522 = notNaN_addZeros & roundingMode_min; // @[MulAddRecFN.scala 291:26:chipyard.TestHarness.RocketConfig.fir@237610.4]
  assign _T_523 = io_fromPreMul_signProd | CDom_sign; // @[MulAddRecFN.scala 292:37:chipyard.TestHarness.RocketConfig.fir@237611.4]
  assign _T_524 = _T_522 & _T_523; // @[MulAddRecFN.scala 291:46:chipyard.TestHarness.RocketConfig.fir@237612.4]
  assign _T_525 = _T_521 | _T_524; // @[MulAddRecFN.scala 290:48:chipyard.TestHarness.RocketConfig.fir@237613.4]
  assign _T_526 = ~notNaN_isInfOut; // @[MulAddRecFN.scala 293:10:chipyard.TestHarness.RocketConfig.fir@237614.4]
  assign _T_527 = ~notNaN_addZeros; // @[MulAddRecFN.scala 293:31:chipyard.TestHarness.RocketConfig.fir@237615.4]
  assign _T_528 = _T_526 & _T_527; // @[MulAddRecFN.scala 293:28:chipyard.TestHarness.RocketConfig.fir@237616.4]
  assign _T_529 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17:chipyard.TestHarness.RocketConfig.fir@237617.4]
  assign _T_530 = _T_528 & _T_529; // @[MulAddRecFN.scala 293:49:chipyard.TestHarness.RocketConfig.fir@237618.4]
  assign io_invalidExc = _T_503 | _T_508; // @[MulAddRecFN.scala 272:19:chipyard.TestHarness.RocketConfig.fir@237594.4]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:21:chipyard.TestHarness.RocketConfig.fir@237596.4]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 281:21:chipyard.TestHarness.RocketConfig.fir@237597.4]
  assign io_rawOut_isZero = notNaN_addZeros | _T_512; // @[MulAddRecFN.scala 283:22:chipyard.TestHarness.RocketConfig.fir@237601.4]
  assign io_rawOut_sign = _T_525 | _T_530; // @[MulAddRecFN.scala 286:20:chipyard.TestHarness.RocketConfig.fir@237620.4]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:20:chipyard.TestHarness.RocketConfig.fir@237622.4]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:19:chipyard.TestHarness.RocketConfig.fir@237624.4]
endmodule
