module MulAddRecFNToRaw_postMul( // @[:chipyard.TestHarness.RocketConfig.fir@233684.2]
  input         io_fromPreMul_isSigNaNAny, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input         io_fromPreMul_isNaNAOrB, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input         io_fromPreMul_isInfA, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input         io_fromPreMul_isZeroA, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input         io_fromPreMul_isInfB, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input         io_fromPreMul_isZeroB, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input         io_fromPreMul_signProd, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input         io_fromPreMul_isNaNC, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input         io_fromPreMul_isInfC, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input         io_fromPreMul_isZeroC, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input  [9:0]  io_fromPreMul_sExpSum, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input         io_fromPreMul_doSubMags, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input         io_fromPreMul_CIsDominant, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input  [4:0]  io_fromPreMul_CDom_CAlignDist, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input  [25:0] io_fromPreMul_highAlignedSigC, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input         io_fromPreMul_bit0AlignedSigC, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input  [48:0] io_mulAddResult, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  input  [2:0]  io_roundingMode, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  output        io_invalidExc, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  output        io_rawOut_isNaN, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  output        io_rawOut_isInf, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  output        io_rawOut_isZero, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  output        io_rawOut_sign, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  output [9:0]  io_rawOut_sExp, // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
  output [26:0] io_rawOut_sig // @[:chipyard.TestHarness.RocketConfig.fir@233685.4]
);
  wire  roundingMode_min; // @[MulAddRecFN.scala 188:45:chipyard.TestHarness.RocketConfig.fir@233688.4]
  wire  CDom_sign; // @[MulAddRecFN.scala 192:42:chipyard.TestHarness.RocketConfig.fir@233689.4]
  wire [25:0] _T_2; // @[MulAddRecFN.scala 195:47:chipyard.TestHarness.RocketConfig.fir@233692.4]
  wire [25:0] _T_3; // @[MulAddRecFN.scala 194:16:chipyard.TestHarness.RocketConfig.fir@233693.4]
  wire [74:0] sigSum; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233696.4]
  wire [1:0] _T_6; // @[MulAddRecFN.scala 205:69:chipyard.TestHarness.RocketConfig.fir@233697.4]
  wire [9:0] _GEN_0; // @[MulAddRecFN.scala 205:43:chipyard.TestHarness.RocketConfig.fir@233698.4]
  wire [9:0] CDom_sExp; // @[MulAddRecFN.scala 205:43:chipyard.TestHarness.RocketConfig.fir@233700.4]
  wire [49:0] _T_10; // @[MulAddRecFN.scala 208:13:chipyard.TestHarness.RocketConfig.fir@233702.4]
  wire [49:0] _T_14; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233706.4]
  wire [49:0] CDom_absSigSum; // @[MulAddRecFN.scala 207:12:chipyard.TestHarness.RocketConfig.fir@233707.4]
  wire [23:0] _T_16; // @[MulAddRecFN.scala 217:14:chipyard.TestHarness.RocketConfig.fir@233709.4]
  wire  _T_17; // @[MulAddRecFN.scala 217:36:chipyard.TestHarness.RocketConfig.fir@233710.4]
  wire  _T_19; // @[MulAddRecFN.scala 218:37:chipyard.TestHarness.RocketConfig.fir@233712.4]
  wire  CDom_absSigSumExtra; // @[MulAddRecFN.scala 216:12:chipyard.TestHarness.RocketConfig.fir@233713.4]
  wire [80:0] _GEN_1; // @[MulAddRecFN.scala 221:24:chipyard.TestHarness.RocketConfig.fir@233714.4]
  wire [80:0] _T_20; // @[MulAddRecFN.scala 221:24:chipyard.TestHarness.RocketConfig.fir@233714.4]
  wire [28:0] CDom_mainSig; // @[MulAddRecFN.scala 221:56:chipyard.TestHarness.RocketConfig.fir@233715.4]
  wire [26:0] _T_22; // @[MulAddRecFN.scala 224:53:chipyard.TestHarness.RocketConfig.fir@233717.4]
  wire  _T_25; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233721.4]
  wire  _T_27; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233724.4]
  wire  _T_29; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233727.4]
  wire  _T_31; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233730.4]
  wire  _T_33; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233733.4]
  wire  _T_35; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233736.4]
  wire  _T_37; // @[primitives.scala 124:57:chipyard.TestHarness.RocketConfig.fir@233739.4]
  wire [6:0] _T_43; // @[primitives.scala 125:20:chipyard.TestHarness.RocketConfig.fir@233746.4]
  wire [2:0] _T_45; // @[primitives.scala 51:21:chipyard.TestHarness.RocketConfig.fir@233748.4]
  wire [8:0] _T_46; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@233749.4]
  wire [5:0] _T_62; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233765.4]
  wire [6:0] _GEN_2; // @[MulAddRecFN.scala 224:72:chipyard.TestHarness.RocketConfig.fir@233766.4]
  wire [6:0] _T_63; // @[MulAddRecFN.scala 224:72:chipyard.TestHarness.RocketConfig.fir@233766.4]
  wire  CDom_reduced4SigExtra; // @[MulAddRecFN.scala 225:73:chipyard.TestHarness.RocketConfig.fir@233767.4]
  wire  _T_66; // @[MulAddRecFN.scala 228:32:chipyard.TestHarness.RocketConfig.fir@233770.4]
  wire  _T_67; // @[MulAddRecFN.scala 228:36:chipyard.TestHarness.RocketConfig.fir@233771.4]
  wire  _T_68; // @[MulAddRecFN.scala 228:61:chipyard.TestHarness.RocketConfig.fir@233772.4]
  wire [26:0] CDom_sig; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233773.4]
  wire  notCDom_signSigSum; // @[MulAddRecFN.scala 234:36:chipyard.TestHarness.RocketConfig.fir@233774.4]
  wire [50:0] _T_70; // @[MulAddRecFN.scala 237:13:chipyard.TestHarness.RocketConfig.fir@233776.4]
  wire [50:0] _GEN_3; // @[MulAddRecFN.scala 238:41:chipyard.TestHarness.RocketConfig.fir@233778.4]
  wire [50:0] _T_73; // @[MulAddRecFN.scala 238:41:chipyard.TestHarness.RocketConfig.fir@233779.4]
  wire [50:0] notCDom_absSigSum; // @[MulAddRecFN.scala 236:12:chipyard.TestHarness.RocketConfig.fir@233780.4]
  wire  _T_76; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233784.4]
  wire  _T_78; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233787.4]
  wire  _T_80; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233790.4]
  wire  _T_82; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233793.4]
  wire  _T_84; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233796.4]
  wire  _T_86; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233799.4]
  wire  _T_88; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233802.4]
  wire  _T_90; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233805.4]
  wire  _T_92; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233808.4]
  wire  _T_94; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233811.4]
  wire  _T_96; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233814.4]
  wire  _T_98; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233817.4]
  wire  _T_100; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233820.4]
  wire  _T_102; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233823.4]
  wire  _T_104; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233826.4]
  wire  _T_106; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233829.4]
  wire  _T_108; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233832.4]
  wire  _T_110; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233835.4]
  wire  _T_112; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233838.4]
  wire  _T_114; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233841.4]
  wire  _T_116; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233844.4]
  wire  _T_118; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233847.4]
  wire  _T_120; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233850.4]
  wire  _T_122; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233853.4]
  wire  _T_124; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233856.4]
  wire  _T_126; // @[primitives.scala 107:57:chipyard.TestHarness.RocketConfig.fir@233859.4]
  wire [5:0] _T_131; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@233865.4]
  wire [12:0] _T_138; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@233872.4]
  wire [5:0] _T_143; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@233877.4]
  wire [25:0] notCDom_reduced2AbsSigSum; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@233885.4]
  wire [4:0] _T_177; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233912.4]
  wire [4:0] _T_178; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233913.4]
  wire [4:0] _T_179; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233914.4]
  wire [4:0] _T_180; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233915.4]
  wire [4:0] _T_181; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233916.4]
  wire [4:0] _T_182; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233917.4]
  wire [4:0] _T_183; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233918.4]
  wire [4:0] _T_184; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233919.4]
  wire [4:0] _T_185; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233920.4]
  wire [4:0] _T_186; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233921.4]
  wire [4:0] _T_187; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233922.4]
  wire [4:0] _T_188; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233923.4]
  wire [4:0] _T_189; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233924.4]
  wire [4:0] _T_190; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233925.4]
  wire [4:0] _T_191; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233926.4]
  wire [4:0] _T_192; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233927.4]
  wire [4:0] _T_193; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233928.4]
  wire [4:0] _T_194; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233929.4]
  wire [4:0] _T_195; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233930.4]
  wire [4:0] _T_196; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233931.4]
  wire [4:0] _T_197; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233932.4]
  wire [4:0] _T_198; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233933.4]
  wire [4:0] _T_199; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233934.4]
  wire [4:0] _T_200; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233935.4]
  wire [4:0] notCDom_normDistReduced2; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233936.4]
  wire [5:0] notCDom_nearNormDist; // @[MulAddRecFN.scala 242:56:chipyard.TestHarness.RocketConfig.fir@233937.4]
  wire [6:0] _T_201; // @[MulAddRecFN.scala 243:69:chipyard.TestHarness.RocketConfig.fir@233938.4]
  wire [9:0] _GEN_4; // @[MulAddRecFN.scala 243:46:chipyard.TestHarness.RocketConfig.fir@233939.4]
  wire [9:0] notCDom_sExp; // @[MulAddRecFN.scala 243:46:chipyard.TestHarness.RocketConfig.fir@233941.4]
  wire [113:0] _GEN_5; // @[MulAddRecFN.scala 245:27:chipyard.TestHarness.RocketConfig.fir@233942.4]
  wire [113:0] _T_204; // @[MulAddRecFN.scala 245:27:chipyard.TestHarness.RocketConfig.fir@233942.4]
  wire [28:0] notCDom_mainSig; // @[MulAddRecFN.scala 245:50:chipyard.TestHarness.RocketConfig.fir@233943.4]
  wire  _T_209; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233949.4]
  wire  _T_211; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233952.4]
  wire  _T_213; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233955.4]
  wire  _T_215; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233958.4]
  wire  _T_217; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233961.4]
  wire  _T_219; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233964.4]
  wire  _T_221; // @[primitives.scala 107:57:chipyard.TestHarness.RocketConfig.fir@233967.4]
  wire [6:0] _T_227; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@233974.4]
  wire [3:0] _T_229; // @[primitives.scala 51:21:chipyard.TestHarness.RocketConfig.fir@233976.4]
  wire [16:0] _T_230; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@233977.4]
  wire [5:0] _T_246; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233993.4]
  wire [6:0] _GEN_6; // @[MulAddRecFN.scala 249:78:chipyard.TestHarness.RocketConfig.fir@233994.4]
  wire [6:0] _T_247; // @[MulAddRecFN.scala 249:78:chipyard.TestHarness.RocketConfig.fir@233994.4]
  wire  notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 251:11:chipyard.TestHarness.RocketConfig.fir@233995.4]
  wire  _T_250; // @[MulAddRecFN.scala 254:35:chipyard.TestHarness.RocketConfig.fir@233998.4]
  wire  _T_251; // @[MulAddRecFN.scala 254:39:chipyard.TestHarness.RocketConfig.fir@233999.4]
  wire [26:0] notCDom_sig; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@234000.4]
  wire  notCDom_completeCancellation; // @[MulAddRecFN.scala 257:50:chipyard.TestHarness.RocketConfig.fir@234002.4]
  wire  _T_253; // @[MulAddRecFN.scala 261:36:chipyard.TestHarness.RocketConfig.fir@234003.4]
  wire  notCDom_sign; // @[MulAddRecFN.scala 259:12:chipyard.TestHarness.RocketConfig.fir@234004.4]
  wire  notNaN_isInfProd; // @[MulAddRecFN.scala 266:49:chipyard.TestHarness.RocketConfig.fir@234005.4]
  wire  notNaN_isInfOut; // @[MulAddRecFN.scala 267:44:chipyard.TestHarness.RocketConfig.fir@234006.4]
  wire  _T_254; // @[MulAddRecFN.scala 269:32:chipyard.TestHarness.RocketConfig.fir@234007.4]
  wire  notNaN_addZeros; // @[MulAddRecFN.scala 269:58:chipyard.TestHarness.RocketConfig.fir@234008.4]
  wire  _T_255; // @[MulAddRecFN.scala 274:31:chipyard.TestHarness.RocketConfig.fir@234009.4]
  wire  _T_256; // @[MulAddRecFN.scala 273:35:chipyard.TestHarness.RocketConfig.fir@234010.4]
  wire  _T_257; // @[MulAddRecFN.scala 275:32:chipyard.TestHarness.RocketConfig.fir@234011.4]
  wire  _T_258; // @[MulAddRecFN.scala 274:57:chipyard.TestHarness.RocketConfig.fir@234012.4]
  wire  _T_259; // @[MulAddRecFN.scala 276:10:chipyard.TestHarness.RocketConfig.fir@234013.4]
  wire  _T_261; // @[MulAddRecFN.scala 276:36:chipyard.TestHarness.RocketConfig.fir@234015.4]
  wire  _T_262; // @[MulAddRecFN.scala 277:61:chipyard.TestHarness.RocketConfig.fir@234016.4]
  wire  _T_263; // @[MulAddRecFN.scala 278:35:chipyard.TestHarness.RocketConfig.fir@234017.4]
  wire  _T_266; // @[MulAddRecFN.scala 285:14:chipyard.TestHarness.RocketConfig.fir@234023.4]
  wire  _T_267; // @[MulAddRecFN.scala 285:42:chipyard.TestHarness.RocketConfig.fir@234024.4]
  wire  _T_269; // @[MulAddRecFN.scala 287:27:chipyard.TestHarness.RocketConfig.fir@234027.4]
  wire  _T_270; // @[MulAddRecFN.scala 288:31:chipyard.TestHarness.RocketConfig.fir@234028.4]
  wire  _T_271; // @[MulAddRecFN.scala 287:54:chipyard.TestHarness.RocketConfig.fir@234029.4]
  wire  _T_272; // @[MulAddRecFN.scala 289:29:chipyard.TestHarness.RocketConfig.fir@234030.4]
  wire  _T_273; // @[MulAddRecFN.scala 289:26:chipyard.TestHarness.RocketConfig.fir@234031.4]
  wire  _T_274; // @[MulAddRecFN.scala 289:48:chipyard.TestHarness.RocketConfig.fir@234032.4]
  wire  _T_275; // @[MulAddRecFN.scala 290:36:chipyard.TestHarness.RocketConfig.fir@234033.4]
  wire  _T_276; // @[MulAddRecFN.scala 288:43:chipyard.TestHarness.RocketConfig.fir@234034.4]
  wire  _T_277; // @[MulAddRecFN.scala 291:26:chipyard.TestHarness.RocketConfig.fir@234035.4]
  wire  _T_278; // @[MulAddRecFN.scala 292:37:chipyard.TestHarness.RocketConfig.fir@234036.4]
  wire  _T_279; // @[MulAddRecFN.scala 291:46:chipyard.TestHarness.RocketConfig.fir@234037.4]
  wire  _T_280; // @[MulAddRecFN.scala 290:48:chipyard.TestHarness.RocketConfig.fir@234038.4]
  wire  _T_281; // @[MulAddRecFN.scala 293:10:chipyard.TestHarness.RocketConfig.fir@234039.4]
  wire  _T_282; // @[MulAddRecFN.scala 293:31:chipyard.TestHarness.RocketConfig.fir@234040.4]
  wire  _T_283; // @[MulAddRecFN.scala 293:28:chipyard.TestHarness.RocketConfig.fir@234041.4]
  wire  _T_284; // @[MulAddRecFN.scala 294:17:chipyard.TestHarness.RocketConfig.fir@234042.4]
  wire  _T_285; // @[MulAddRecFN.scala 293:49:chipyard.TestHarness.RocketConfig.fir@234043.4]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[MulAddRecFN.scala 188:45:chipyard.TestHarness.RocketConfig.fir@233688.4]
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42:chipyard.TestHarness.RocketConfig.fir@233689.4]
  assign _T_2 = io_fromPreMul_highAlignedSigC + 26'h1; // @[MulAddRecFN.scala 195:47:chipyard.TestHarness.RocketConfig.fir@233692.4]
  assign _T_3 = io_mulAddResult[48] ? _T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16:chipyard.TestHarness.RocketConfig.fir@233693.4]
  assign sigSum = {_T_3,io_mulAddResult[47:0],io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233696.4]
  assign _T_6 = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69:chipyard.TestHarness.RocketConfig.fir@233697.4]
  assign _GEN_0 = {{8{_T_6[1]}},_T_6}; // @[MulAddRecFN.scala 205:43:chipyard.TestHarness.RocketConfig.fir@233698.4]
  assign CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43:chipyard.TestHarness.RocketConfig.fir@233700.4]
  assign _T_10 = ~sigSum[74:25]; // @[MulAddRecFN.scala 208:13:chipyard.TestHarness.RocketConfig.fir@233702.4]
  assign _T_14 = {1'h0,io_fromPreMul_highAlignedSigC[25:24],sigSum[72:26]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233706.4]
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? _T_10 : _T_14; // @[MulAddRecFN.scala 207:12:chipyard.TestHarness.RocketConfig.fir@233707.4]
  assign _T_16 = ~sigSum[24:1]; // @[MulAddRecFN.scala 217:14:chipyard.TestHarness.RocketConfig.fir@233709.4]
  assign _T_17 = |_T_16; // @[MulAddRecFN.scala 217:36:chipyard.TestHarness.RocketConfig.fir@233710.4]
  assign _T_19 = |sigSum[25:1]; // @[MulAddRecFN.scala 218:37:chipyard.TestHarness.RocketConfig.fir@233712.4]
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _T_17 : _T_19; // @[MulAddRecFN.scala 216:12:chipyard.TestHarness.RocketConfig.fir@233713.4]
  assign _GEN_1 = {{31'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24:chipyard.TestHarness.RocketConfig.fir@233714.4]
  assign _T_20 = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24:chipyard.TestHarness.RocketConfig.fir@233714.4]
  assign CDom_mainSig = _T_20[49:21]; // @[MulAddRecFN.scala 221:56:chipyard.TestHarness.RocketConfig.fir@233715.4]
  assign _T_22 = {CDom_absSigSum[23:0], 3'h0}; // @[MulAddRecFN.scala 224:53:chipyard.TestHarness.RocketConfig.fir@233717.4]
  assign _T_25 = |_T_22[3:0]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233721.4]
  assign _T_27 = |_T_22[7:4]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233724.4]
  assign _T_29 = |_T_22[11:8]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233727.4]
  assign _T_31 = |_T_22[15:12]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233730.4]
  assign _T_33 = |_T_22[19:16]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233733.4]
  assign _T_35 = |_T_22[23:20]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233736.4]
  assign _T_37 = |_T_22[26:24]; // @[primitives.scala 124:57:chipyard.TestHarness.RocketConfig.fir@233739.4]
  assign _T_43 = {_T_37,_T_35,_T_33,_T_31,_T_29,_T_27,_T_25}; // @[primitives.scala 125:20:chipyard.TestHarness.RocketConfig.fir@233746.4]
  assign _T_45 = ~io_fromPreMul_CDom_CAlignDist[4:2]; // @[primitives.scala 51:21:chipyard.TestHarness.RocketConfig.fir@233748.4]
  assign _T_46 = -9'sh100 >>> _T_45; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@233749.4]
  assign _T_62 = {_T_46[1],_T_46[2],_T_46[3],_T_46[4],_T_46[5],_T_46[6]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233765.4]
  assign _GEN_2 = {{1'd0}, _T_62}; // @[MulAddRecFN.scala 224:72:chipyard.TestHarness.RocketConfig.fir@233766.4]
  assign _T_63 = _T_43 & _GEN_2; // @[MulAddRecFN.scala 224:72:chipyard.TestHarness.RocketConfig.fir@233766.4]
  assign CDom_reduced4SigExtra = |_T_63; // @[MulAddRecFN.scala 225:73:chipyard.TestHarness.RocketConfig.fir@233767.4]
  assign _T_66 = |CDom_mainSig[2:0]; // @[MulAddRecFN.scala 228:32:chipyard.TestHarness.RocketConfig.fir@233770.4]
  assign _T_67 = _T_66 | CDom_reduced4SigExtra; // @[MulAddRecFN.scala 228:36:chipyard.TestHarness.RocketConfig.fir@233771.4]
  assign _T_68 = _T_67 | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61:chipyard.TestHarness.RocketConfig.fir@233772.4]
  assign CDom_sig = {CDom_mainSig[28:3],_T_68}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233773.4]
  assign notCDom_signSigSum = sigSum[51]; // @[MulAddRecFN.scala 234:36:chipyard.TestHarness.RocketConfig.fir@233774.4]
  assign _T_70 = ~sigSum[50:0]; // @[MulAddRecFN.scala 237:13:chipyard.TestHarness.RocketConfig.fir@233776.4]
  assign _GEN_3 = {{50'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41:chipyard.TestHarness.RocketConfig.fir@233778.4]
  assign _T_73 = sigSum[50:0] + _GEN_3; // @[MulAddRecFN.scala 238:41:chipyard.TestHarness.RocketConfig.fir@233779.4]
  assign notCDom_absSigSum = notCDom_signSigSum ? _T_70 : _T_73; // @[MulAddRecFN.scala 236:12:chipyard.TestHarness.RocketConfig.fir@233780.4]
  assign _T_76 = |notCDom_absSigSum[1:0]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233784.4]
  assign _T_78 = |notCDom_absSigSum[3:2]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233787.4]
  assign _T_80 = |notCDom_absSigSum[5:4]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233790.4]
  assign _T_82 = |notCDom_absSigSum[7:6]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233793.4]
  assign _T_84 = |notCDom_absSigSum[9:8]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233796.4]
  assign _T_86 = |notCDom_absSigSum[11:10]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233799.4]
  assign _T_88 = |notCDom_absSigSum[13:12]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233802.4]
  assign _T_90 = |notCDom_absSigSum[15:14]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233805.4]
  assign _T_92 = |notCDom_absSigSum[17:16]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233808.4]
  assign _T_94 = |notCDom_absSigSum[19:18]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233811.4]
  assign _T_96 = |notCDom_absSigSum[21:20]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233814.4]
  assign _T_98 = |notCDom_absSigSum[23:22]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233817.4]
  assign _T_100 = |notCDom_absSigSum[25:24]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233820.4]
  assign _T_102 = |notCDom_absSigSum[27:26]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233823.4]
  assign _T_104 = |notCDom_absSigSum[29:28]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233826.4]
  assign _T_106 = |notCDom_absSigSum[31:30]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233829.4]
  assign _T_108 = |notCDom_absSigSum[33:32]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233832.4]
  assign _T_110 = |notCDom_absSigSum[35:34]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233835.4]
  assign _T_112 = |notCDom_absSigSum[37:36]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233838.4]
  assign _T_114 = |notCDom_absSigSum[39:38]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233841.4]
  assign _T_116 = |notCDom_absSigSum[41:40]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233844.4]
  assign _T_118 = |notCDom_absSigSum[43:42]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233847.4]
  assign _T_120 = |notCDom_absSigSum[45:44]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233850.4]
  assign _T_122 = |notCDom_absSigSum[47:46]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233853.4]
  assign _T_124 = |notCDom_absSigSum[49:48]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233856.4]
  assign _T_126 = |notCDom_absSigSum[50]; // @[primitives.scala 107:57:chipyard.TestHarness.RocketConfig.fir@233859.4]
  assign _T_131 = {_T_86,_T_84,_T_82,_T_80,_T_78,_T_76}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@233865.4]
  assign _T_138 = {_T_100,_T_98,_T_96,_T_94,_T_92,_T_90,_T_88,_T_131}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@233872.4]
  assign _T_143 = {_T_112,_T_110,_T_108,_T_106,_T_104,_T_102}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@233877.4]
  assign notCDom_reduced2AbsSigSum = {_T_126,_T_124,_T_122,_T_120,_T_118,_T_116,_T_114,_T_143,_T_138}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@233885.4]
  assign _T_177 = notCDom_reduced2AbsSigSum[1] ? 5'h18 : 5'h19; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233912.4]
  assign _T_178 = notCDom_reduced2AbsSigSum[2] ? 5'h17 : _T_177; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233913.4]
  assign _T_179 = notCDom_reduced2AbsSigSum[3] ? 5'h16 : _T_178; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233914.4]
  assign _T_180 = notCDom_reduced2AbsSigSum[4] ? 5'h15 : _T_179; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233915.4]
  assign _T_181 = notCDom_reduced2AbsSigSum[5] ? 5'h14 : _T_180; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233916.4]
  assign _T_182 = notCDom_reduced2AbsSigSum[6] ? 5'h13 : _T_181; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233917.4]
  assign _T_183 = notCDom_reduced2AbsSigSum[7] ? 5'h12 : _T_182; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233918.4]
  assign _T_184 = notCDom_reduced2AbsSigSum[8] ? 5'h11 : _T_183; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233919.4]
  assign _T_185 = notCDom_reduced2AbsSigSum[9] ? 5'h10 : _T_184; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233920.4]
  assign _T_186 = notCDom_reduced2AbsSigSum[10] ? 5'hf : _T_185; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233921.4]
  assign _T_187 = notCDom_reduced2AbsSigSum[11] ? 5'he : _T_186; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233922.4]
  assign _T_188 = notCDom_reduced2AbsSigSum[12] ? 5'hd : _T_187; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233923.4]
  assign _T_189 = notCDom_reduced2AbsSigSum[13] ? 5'hc : _T_188; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233924.4]
  assign _T_190 = notCDom_reduced2AbsSigSum[14] ? 5'hb : _T_189; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233925.4]
  assign _T_191 = notCDom_reduced2AbsSigSum[15] ? 5'ha : _T_190; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233926.4]
  assign _T_192 = notCDom_reduced2AbsSigSum[16] ? 5'h9 : _T_191; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233927.4]
  assign _T_193 = notCDom_reduced2AbsSigSum[17] ? 5'h8 : _T_192; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233928.4]
  assign _T_194 = notCDom_reduced2AbsSigSum[18] ? 5'h7 : _T_193; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233929.4]
  assign _T_195 = notCDom_reduced2AbsSigSum[19] ? 5'h6 : _T_194; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233930.4]
  assign _T_196 = notCDom_reduced2AbsSigSum[20] ? 5'h5 : _T_195; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233931.4]
  assign _T_197 = notCDom_reduced2AbsSigSum[21] ? 5'h4 : _T_196; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233932.4]
  assign _T_198 = notCDom_reduced2AbsSigSum[22] ? 5'h3 : _T_197; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233933.4]
  assign _T_199 = notCDom_reduced2AbsSigSum[23] ? 5'h2 : _T_198; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233934.4]
  assign _T_200 = notCDom_reduced2AbsSigSum[24] ? 5'h1 : _T_199; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233935.4]
  assign notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[25] ? 5'h0 : _T_200; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@233936.4]
  assign notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56:chipyard.TestHarness.RocketConfig.fir@233937.4]
  assign _T_201 = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69:chipyard.TestHarness.RocketConfig.fir@233938.4]
  assign _GEN_4 = {{3{_T_201[6]}},_T_201}; // @[MulAddRecFN.scala 243:46:chipyard.TestHarness.RocketConfig.fir@233939.4]
  assign notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_4); // @[MulAddRecFN.scala 243:46:chipyard.TestHarness.RocketConfig.fir@233941.4]
  assign _GEN_5 = {{63'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27:chipyard.TestHarness.RocketConfig.fir@233942.4]
  assign _T_204 = _GEN_5 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27:chipyard.TestHarness.RocketConfig.fir@233942.4]
  assign notCDom_mainSig = _T_204[51:23]; // @[MulAddRecFN.scala 245:50:chipyard.TestHarness.RocketConfig.fir@233943.4]
  assign _T_209 = |notCDom_reduced2AbsSigSum[1:0]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233949.4]
  assign _T_211 = |notCDom_reduced2AbsSigSum[3:2]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233952.4]
  assign _T_213 = |notCDom_reduced2AbsSigSum[5:4]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233955.4]
  assign _T_215 = |notCDom_reduced2AbsSigSum[7:6]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233958.4]
  assign _T_217 = |notCDom_reduced2AbsSigSum[9:8]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233961.4]
  assign _T_219 = |notCDom_reduced2AbsSigSum[11:10]; // @[primitives.scala 104:54:chipyard.TestHarness.RocketConfig.fir@233964.4]
  assign _T_221 = |notCDom_reduced2AbsSigSum[12]; // @[primitives.scala 107:57:chipyard.TestHarness.RocketConfig.fir@233967.4]
  assign _T_227 = {_T_221,_T_219,_T_217,_T_215,_T_213,_T_211,_T_209}; // @[primitives.scala 108:20:chipyard.TestHarness.RocketConfig.fir@233974.4]
  assign _T_229 = ~notCDom_normDistReduced2[4:1]; // @[primitives.scala 51:21:chipyard.TestHarness.RocketConfig.fir@233976.4]
  assign _T_230 = -17'sh10000 >>> _T_229; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@233977.4]
  assign _T_246 = {_T_230[1],_T_230[2],_T_230[3],_T_230[4],_T_230[5],_T_230[6]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233993.4]
  assign _GEN_6 = {{1'd0}, _T_246}; // @[MulAddRecFN.scala 249:78:chipyard.TestHarness.RocketConfig.fir@233994.4]
  assign _T_247 = _T_227 & _GEN_6; // @[MulAddRecFN.scala 249:78:chipyard.TestHarness.RocketConfig.fir@233994.4]
  assign notCDom_reduced4SigExtra = |_T_247; // @[MulAddRecFN.scala 251:11:chipyard.TestHarness.RocketConfig.fir@233995.4]
  assign _T_250 = |notCDom_mainSig[2:0]; // @[MulAddRecFN.scala 254:35:chipyard.TestHarness.RocketConfig.fir@233998.4]
  assign _T_251 = _T_250 | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39:chipyard.TestHarness.RocketConfig.fir@233999.4]
  assign notCDom_sig = {notCDom_mainSig[28:3],_T_251}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@234000.4]
  assign notCDom_completeCancellation = notCDom_sig[26:25] == 2'h0; // @[MulAddRecFN.scala 257:50:chipyard.TestHarness.RocketConfig.fir@234002.4]
  assign _T_253 = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36:chipyard.TestHarness.RocketConfig.fir@234003.4]
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : _T_253; // @[MulAddRecFN.scala 259:12:chipyard.TestHarness.RocketConfig.fir@234004.4]
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49:chipyard.TestHarness.RocketConfig.fir@234005.4]
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44:chipyard.TestHarness.RocketConfig.fir@234006.4]
  assign _T_254 = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 269:32:chipyard.TestHarness.RocketConfig.fir@234007.4]
  assign notNaN_addZeros = _T_254 & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58:chipyard.TestHarness.RocketConfig.fir@234008.4]
  assign _T_255 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31:chipyard.TestHarness.RocketConfig.fir@234009.4]
  assign _T_256 = io_fromPreMul_isSigNaNAny | _T_255; // @[MulAddRecFN.scala 273:35:chipyard.TestHarness.RocketConfig.fir@234010.4]
  assign _T_257 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32:chipyard.TestHarness.RocketConfig.fir@234011.4]
  assign _T_258 = _T_256 | _T_257; // @[MulAddRecFN.scala 274:57:chipyard.TestHarness.RocketConfig.fir@234012.4]
  assign _T_259 = ~io_fromPreMul_isNaNAOrB; // @[MulAddRecFN.scala 276:10:chipyard.TestHarness.RocketConfig.fir@234013.4]
  assign _T_261 = _T_259 & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36:chipyard.TestHarness.RocketConfig.fir@234015.4]
  assign _T_262 = _T_261 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61:chipyard.TestHarness.RocketConfig.fir@234016.4]
  assign _T_263 = _T_262 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35:chipyard.TestHarness.RocketConfig.fir@234017.4]
  assign _T_266 = ~io_fromPreMul_CIsDominant; // @[MulAddRecFN.scala 285:14:chipyard.TestHarness.RocketConfig.fir@234023.4]
  assign _T_267 = _T_266 & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42:chipyard.TestHarness.RocketConfig.fir@234024.4]
  assign _T_269 = notNaN_isInfProd & io_fromPreMul_signProd; // @[MulAddRecFN.scala 287:27:chipyard.TestHarness.RocketConfig.fir@234027.4]
  assign _T_270 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31:chipyard.TestHarness.RocketConfig.fir@234028.4]
  assign _T_271 = _T_269 | _T_270; // @[MulAddRecFN.scala 287:54:chipyard.TestHarness.RocketConfig.fir@234029.4]
  assign _T_272 = ~roundingMode_min; // @[MulAddRecFN.scala 289:29:chipyard.TestHarness.RocketConfig.fir@234030.4]
  assign _T_273 = notNaN_addZeros & _T_272; // @[MulAddRecFN.scala 289:26:chipyard.TestHarness.RocketConfig.fir@234031.4]
  assign _T_274 = _T_273 & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48:chipyard.TestHarness.RocketConfig.fir@234032.4]
  assign _T_275 = _T_274 & CDom_sign; // @[MulAddRecFN.scala 290:36:chipyard.TestHarness.RocketConfig.fir@234033.4]
  assign _T_276 = _T_271 | _T_275; // @[MulAddRecFN.scala 288:43:chipyard.TestHarness.RocketConfig.fir@234034.4]
  assign _T_277 = notNaN_addZeros & roundingMode_min; // @[MulAddRecFN.scala 291:26:chipyard.TestHarness.RocketConfig.fir@234035.4]
  assign _T_278 = io_fromPreMul_signProd | CDom_sign; // @[MulAddRecFN.scala 292:37:chipyard.TestHarness.RocketConfig.fir@234036.4]
  assign _T_279 = _T_277 & _T_278; // @[MulAddRecFN.scala 291:46:chipyard.TestHarness.RocketConfig.fir@234037.4]
  assign _T_280 = _T_276 | _T_279; // @[MulAddRecFN.scala 290:48:chipyard.TestHarness.RocketConfig.fir@234038.4]
  assign _T_281 = ~notNaN_isInfOut; // @[MulAddRecFN.scala 293:10:chipyard.TestHarness.RocketConfig.fir@234039.4]
  assign _T_282 = ~notNaN_addZeros; // @[MulAddRecFN.scala 293:31:chipyard.TestHarness.RocketConfig.fir@234040.4]
  assign _T_283 = _T_281 & _T_282; // @[MulAddRecFN.scala 293:28:chipyard.TestHarness.RocketConfig.fir@234041.4]
  assign _T_284 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17:chipyard.TestHarness.RocketConfig.fir@234042.4]
  assign _T_285 = _T_283 & _T_284; // @[MulAddRecFN.scala 293:49:chipyard.TestHarness.RocketConfig.fir@234043.4]
  assign io_invalidExc = _T_258 | _T_263; // @[MulAddRecFN.scala 272:19:chipyard.TestHarness.RocketConfig.fir@234019.4]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:21:chipyard.TestHarness.RocketConfig.fir@234021.4]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 281:21:chipyard.TestHarness.RocketConfig.fir@234022.4]
  assign io_rawOut_isZero = notNaN_addZeros | _T_267; // @[MulAddRecFN.scala 283:22:chipyard.TestHarness.RocketConfig.fir@234026.4]
  assign io_rawOut_sign = _T_280 | _T_285; // @[MulAddRecFN.scala 286:20:chipyard.TestHarness.RocketConfig.fir@234045.4]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:20:chipyard.TestHarness.RocketConfig.fir@234047.4]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:19:chipyard.TestHarness.RocketConfig.fir@234049.4]
endmodule
