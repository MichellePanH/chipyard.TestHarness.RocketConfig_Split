module MulAddRecFNToRaw_preMul( // @[:chipyard.TestHarness.RocketConfig.fir@233475.2]
  input  [1:0]  io_op, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  input  [32:0] io_a, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  input  [32:0] io_b, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  input  [32:0] io_c, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output [23:0] io_mulAddA, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output [23:0] io_mulAddB, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output [47:0] io_mulAddC, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output        io_toPostMul_isSigNaNAny, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output        io_toPostMul_isNaNAOrB, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output        io_toPostMul_isInfA, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output        io_toPostMul_isZeroA, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output        io_toPostMul_isInfB, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output        io_toPostMul_isZeroB, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output        io_toPostMul_signProd, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output        io_toPostMul_isNaNC, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output        io_toPostMul_isInfC, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output        io_toPostMul_isZeroC, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output [9:0]  io_toPostMul_sExpSum, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output        io_toPostMul_doSubMags, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output        io_toPostMul_CIsDominant, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output [4:0]  io_toPostMul_CDom_CAlignDist, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output [25:0] io_toPostMul_highAlignedSigC, // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
  output        io_toPostMul_bit0AlignedSigC // @[:chipyard.TestHarness.RocketConfig.fir@233476.4]
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54:chipyard.TestHarness.RocketConfig.fir@233481.4]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54:chipyard.TestHarness.RocketConfig.fir@233483.4]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33:chipyard.TestHarness.RocketConfig.fir@233487.4]
  wire  _T_8; // @[rawFloatFromRecFN.scala 56:36:chipyard.TestHarness.RocketConfig.fir@233490.4]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25:chipyard.TestHarness.RocketConfig.fir@233494.4]
  wire [9:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27:chipyard.TestHarness.RocketConfig.fir@233496.4]
  wire  _T_12; // @[rawFloatFromRecFN.scala 60:39:chipyard.TestHarness.RocketConfig.fir@233498.4]
  wire [24:0] rawA_sig; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233501.4]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54:chipyard.TestHarness.RocketConfig.fir@233505.4]
  wire  _T_20; // @[rawFloatFromRecFN.scala 52:54:chipyard.TestHarness.RocketConfig.fir@233507.4]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33:chipyard.TestHarness.RocketConfig.fir@233511.4]
  wire  _T_24; // @[rawFloatFromRecFN.scala 56:36:chipyard.TestHarness.RocketConfig.fir@233514.4]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25:chipyard.TestHarness.RocketConfig.fir@233518.4]
  wire [9:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27:chipyard.TestHarness.RocketConfig.fir@233520.4]
  wire  _T_28; // @[rawFloatFromRecFN.scala 60:39:chipyard.TestHarness.RocketConfig.fir@233522.4]
  wire [24:0] rawB_sig; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233525.4]
  wire  rawC_isZero; // @[rawFloatFromRecFN.scala 51:54:chipyard.TestHarness.RocketConfig.fir@233529.4]
  wire  _T_36; // @[rawFloatFromRecFN.scala 52:54:chipyard.TestHarness.RocketConfig.fir@233531.4]
  wire  rawC_isNaN; // @[rawFloatFromRecFN.scala 55:33:chipyard.TestHarness.RocketConfig.fir@233535.4]
  wire  _T_40; // @[rawFloatFromRecFN.scala 56:36:chipyard.TestHarness.RocketConfig.fir@233538.4]
  wire  rawC_sign; // @[rawFloatFromRecFN.scala 58:25:chipyard.TestHarness.RocketConfig.fir@233542.4]
  wire [9:0] rawC_sExp; // @[rawFloatFromRecFN.scala 59:27:chipyard.TestHarness.RocketConfig.fir@233544.4]
  wire  _T_44; // @[rawFloatFromRecFN.scala 60:39:chipyard.TestHarness.RocketConfig.fir@233546.4]
  wire [24:0] rawC_sig; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233549.4]
  wire  _T_48; // @[MulAddRecFN.scala 98:30:chipyard.TestHarness.RocketConfig.fir@233551.4]
  wire  signProd; // @[MulAddRecFN.scala 98:42:chipyard.TestHarness.RocketConfig.fir@233553.4]
  wire [10:0] _T_50; // @[MulAddRecFN.scala 101:19:chipyard.TestHarness.RocketConfig.fir@233554.4]
  wire [10:0] sExpAlignedProd; // @[MulAddRecFN.scala 101:32:chipyard.TestHarness.RocketConfig.fir@233557.4]
  wire  _T_53; // @[MulAddRecFN.scala 103:30:chipyard.TestHarness.RocketConfig.fir@233558.4]
  wire  doSubMags; // @[MulAddRecFN.scala 103:42:chipyard.TestHarness.RocketConfig.fir@233560.4]
  wire [10:0] _GEN_0; // @[MulAddRecFN.scala 107:42:chipyard.TestHarness.RocketConfig.fir@233561.4]
  wire [10:0] sNatCAlignDist; // @[MulAddRecFN.scala 107:42:chipyard.TestHarness.RocketConfig.fir@233563.4]
  wire [9:0] posNatCAlignDist; // @[MulAddRecFN.scala 108:42:chipyard.TestHarness.RocketConfig.fir@233564.4]
  wire  _T_57; // @[MulAddRecFN.scala 109:35:chipyard.TestHarness.RocketConfig.fir@233565.4]
  wire  _T_58; // @[MulAddRecFN.scala 109:69:chipyard.TestHarness.RocketConfig.fir@233566.4]
  wire  isMinCAlign; // @[MulAddRecFN.scala 109:50:chipyard.TestHarness.RocketConfig.fir@233567.4]
  wire  _T_60; // @[MulAddRecFN.scala 111:60:chipyard.TestHarness.RocketConfig.fir@233569.4]
  wire  _T_61; // @[MulAddRecFN.scala 111:39:chipyard.TestHarness.RocketConfig.fir@233570.4]
  wire  CIsDominant; // @[MulAddRecFN.scala 111:23:chipyard.TestHarness.RocketConfig.fir@233571.4]
  wire  _T_62; // @[MulAddRecFN.scala 115:34:chipyard.TestHarness.RocketConfig.fir@233572.4]
  wire [6:0] _T_64; // @[MulAddRecFN.scala 115:16:chipyard.TestHarness.RocketConfig.fir@233574.4]
  wire [6:0] CAlignDist; // @[MulAddRecFN.scala 113:12:chipyard.TestHarness.RocketConfig.fir@233575.4]
  wire [24:0] _T_65; // @[MulAddRecFN.scala 121:28:chipyard.TestHarness.RocketConfig.fir@233576.4]
  wire [24:0] _T_66; // @[MulAddRecFN.scala 121:16:chipyard.TestHarness.RocketConfig.fir@233577.4]
  wire [52:0] _T_68; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@233579.4]
  wire [77:0] _T_70; // @[MulAddRecFN.scala 123:11:chipyard.TestHarness.RocketConfig.fir@233581.4]
  wire [77:0] mainAlignedSigC; // @[MulAddRecFN.scala 123:17:chipyard.TestHarness.RocketConfig.fir@233582.4]
  wire [26:0] _T_71; // @[MulAddRecFN.scala 125:30:chipyard.TestHarness.RocketConfig.fir@233583.4]
  wire  _T_74; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233587.4]
  wire  _T_76; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233590.4]
  wire  _T_78; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233593.4]
  wire  _T_80; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233596.4]
  wire  _T_82; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233599.4]
  wire  _T_84; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233602.4]
  wire  _T_86; // @[primitives.scala 124:57:chipyard.TestHarness.RocketConfig.fir@233605.4]
  wire [6:0] _T_92; // @[primitives.scala 125:20:chipyard.TestHarness.RocketConfig.fir@233612.4]
  wire [32:0] _T_94; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@233614.4]
  wire [5:0] _T_110; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233630.4]
  wire [6:0] _GEN_1; // @[MulAddRecFN.scala 125:68:chipyard.TestHarness.RocketConfig.fir@233631.4]
  wire [6:0] _T_111; // @[MulAddRecFN.scala 125:68:chipyard.TestHarness.RocketConfig.fir@233631.4]
  wire  reduced4CExtra; // @[MulAddRecFN.scala 133:11:chipyard.TestHarness.RocketConfig.fir@233632.4]
  wire  _T_114; // @[MulAddRecFN.scala 137:39:chipyard.TestHarness.RocketConfig.fir@233635.4]
  wire  _T_115; // @[MulAddRecFN.scala 137:47:chipyard.TestHarness.RocketConfig.fir@233636.4]
  wire  _T_116; // @[MulAddRecFN.scala 137:44:chipyard.TestHarness.RocketConfig.fir@233637.4]
  wire  _T_118; // @[MulAddRecFN.scala 138:39:chipyard.TestHarness.RocketConfig.fir@233639.4]
  wire  _T_119; // @[MulAddRecFN.scala 138:44:chipyard.TestHarness.RocketConfig.fir@233640.4]
  wire  _T_120; // @[MulAddRecFN.scala 136:16:chipyard.TestHarness.RocketConfig.fir@233641.4]
  wire [74:0] _T_121; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233642.4]
  wire [75:0] alignedSigC; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233643.4]
  wire  _T_124; // @[common.scala 81:49:chipyard.TestHarness.RocketConfig.fir@233649.4]
  wire  _T_125; // @[common.scala 81:46:chipyard.TestHarness.RocketConfig.fir@233650.4]
  wire  _T_127; // @[common.scala 81:49:chipyard.TestHarness.RocketConfig.fir@233652.4]
  wire  _T_128; // @[common.scala 81:46:chipyard.TestHarness.RocketConfig.fir@233653.4]
  wire  _T_129; // @[MulAddRecFN.scala 149:32:chipyard.TestHarness.RocketConfig.fir@233654.4]
  wire  _T_131; // @[common.scala 81:49:chipyard.TestHarness.RocketConfig.fir@233656.4]
  wire  _T_132; // @[common.scala 81:46:chipyard.TestHarness.RocketConfig.fir@233657.4]
  wire [10:0] _T_137; // @[MulAddRecFN.scala 161:53:chipyard.TestHarness.RocketConfig.fir@233672.4]
  wire [10:0] _T_138; // @[MulAddRecFN.scala 161:12:chipyard.TestHarness.RocketConfig.fir@233673.4]
  assign rawA_isZero = io_a[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54:chipyard.TestHarness.RocketConfig.fir@233481.4]
  assign _T_4 = io_a[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54:chipyard.TestHarness.RocketConfig.fir@233483.4]
  assign rawA_isNaN = _T_4 & io_a[29]; // @[rawFloatFromRecFN.scala 55:33:chipyard.TestHarness.RocketConfig.fir@233487.4]
  assign _T_8 = ~io_a[29]; // @[rawFloatFromRecFN.scala 56:36:chipyard.TestHarness.RocketConfig.fir@233490.4]
  assign rawA_sign = io_a[32]; // @[rawFloatFromRecFN.scala 58:25:chipyard.TestHarness.RocketConfig.fir@233494.4]
  assign rawA_sExp = {1'b0,$signed(io_a[31:23])}; // @[rawFloatFromRecFN.scala 59:27:chipyard.TestHarness.RocketConfig.fir@233496.4]
  assign _T_12 = ~rawA_isZero; // @[rawFloatFromRecFN.scala 60:39:chipyard.TestHarness.RocketConfig.fir@233498.4]
  assign rawA_sig = {1'h0,_T_12,io_a[22:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233501.4]
  assign rawB_isZero = io_b[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54:chipyard.TestHarness.RocketConfig.fir@233505.4]
  assign _T_20 = io_b[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54:chipyard.TestHarness.RocketConfig.fir@233507.4]
  assign rawB_isNaN = _T_20 & io_b[29]; // @[rawFloatFromRecFN.scala 55:33:chipyard.TestHarness.RocketConfig.fir@233511.4]
  assign _T_24 = ~io_b[29]; // @[rawFloatFromRecFN.scala 56:36:chipyard.TestHarness.RocketConfig.fir@233514.4]
  assign rawB_sign = io_b[32]; // @[rawFloatFromRecFN.scala 58:25:chipyard.TestHarness.RocketConfig.fir@233518.4]
  assign rawB_sExp = {1'b0,$signed(io_b[31:23])}; // @[rawFloatFromRecFN.scala 59:27:chipyard.TestHarness.RocketConfig.fir@233520.4]
  assign _T_28 = ~rawB_isZero; // @[rawFloatFromRecFN.scala 60:39:chipyard.TestHarness.RocketConfig.fir@233522.4]
  assign rawB_sig = {1'h0,_T_28,io_b[22:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233525.4]
  assign rawC_isZero = io_c[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54:chipyard.TestHarness.RocketConfig.fir@233529.4]
  assign _T_36 = io_c[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54:chipyard.TestHarness.RocketConfig.fir@233531.4]
  assign rawC_isNaN = _T_36 & io_c[29]; // @[rawFloatFromRecFN.scala 55:33:chipyard.TestHarness.RocketConfig.fir@233535.4]
  assign _T_40 = ~io_c[29]; // @[rawFloatFromRecFN.scala 56:36:chipyard.TestHarness.RocketConfig.fir@233538.4]
  assign rawC_sign = io_c[32]; // @[rawFloatFromRecFN.scala 58:25:chipyard.TestHarness.RocketConfig.fir@233542.4]
  assign rawC_sExp = {1'b0,$signed(io_c[31:23])}; // @[rawFloatFromRecFN.scala 59:27:chipyard.TestHarness.RocketConfig.fir@233544.4]
  assign _T_44 = ~rawC_isZero; // @[rawFloatFromRecFN.scala 60:39:chipyard.TestHarness.RocketConfig.fir@233546.4]
  assign rawC_sig = {1'h0,_T_44,io_c[22:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233549.4]
  assign _T_48 = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30:chipyard.TestHarness.RocketConfig.fir@233551.4]
  assign signProd = _T_48 ^ io_op[1]; // @[MulAddRecFN.scala 98:42:chipyard.TestHarness.RocketConfig.fir@233553.4]
  assign _T_50 = $signed(rawA_sExp) + $signed(rawB_sExp); // @[MulAddRecFN.scala 101:19:chipyard.TestHarness.RocketConfig.fir@233554.4]
  assign sExpAlignedProd = $signed(_T_50) - 11'she5; // @[MulAddRecFN.scala 101:32:chipyard.TestHarness.RocketConfig.fir@233557.4]
  assign _T_53 = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30:chipyard.TestHarness.RocketConfig.fir@233558.4]
  assign doSubMags = _T_53 ^ io_op[0]; // @[MulAddRecFN.scala 103:42:chipyard.TestHarness.RocketConfig.fir@233560.4]
  assign _GEN_0 = {{1{rawC_sExp[9]}},rawC_sExp}; // @[MulAddRecFN.scala 107:42:chipyard.TestHarness.RocketConfig.fir@233561.4]
  assign sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42:chipyard.TestHarness.RocketConfig.fir@233563.4]
  assign posNatCAlignDist = sNatCAlignDist[9:0]; // @[MulAddRecFN.scala 108:42:chipyard.TestHarness.RocketConfig.fir@233564.4]
  assign _T_57 = rawA_isZero | rawB_isZero; // @[MulAddRecFN.scala 109:35:chipyard.TestHarness.RocketConfig.fir@233565.4]
  assign _T_58 = $signed(sNatCAlignDist) < 11'sh0; // @[MulAddRecFN.scala 109:69:chipyard.TestHarness.RocketConfig.fir@233566.4]
  assign isMinCAlign = _T_57 | _T_58; // @[MulAddRecFN.scala 109:50:chipyard.TestHarness.RocketConfig.fir@233567.4]
  assign _T_60 = posNatCAlignDist <= 10'h18; // @[MulAddRecFN.scala 111:60:chipyard.TestHarness.RocketConfig.fir@233569.4]
  assign _T_61 = isMinCAlign | _T_60; // @[MulAddRecFN.scala 111:39:chipyard.TestHarness.RocketConfig.fir@233570.4]
  assign CIsDominant = _T_44 & _T_61; // @[MulAddRecFN.scala 111:23:chipyard.TestHarness.RocketConfig.fir@233571.4]
  assign _T_62 = posNatCAlignDist < 10'h4a; // @[MulAddRecFN.scala 115:34:chipyard.TestHarness.RocketConfig.fir@233572.4]
  assign _T_64 = _T_62 ? posNatCAlignDist[6:0] : 7'h4a; // @[MulAddRecFN.scala 115:16:chipyard.TestHarness.RocketConfig.fir@233574.4]
  assign CAlignDist = isMinCAlign ? 7'h0 : _T_64; // @[MulAddRecFN.scala 113:12:chipyard.TestHarness.RocketConfig.fir@233575.4]
  assign _T_65 = ~rawC_sig; // @[MulAddRecFN.scala 121:28:chipyard.TestHarness.RocketConfig.fir@233576.4]
  assign _T_66 = doSubMags ? _T_65 : rawC_sig; // @[MulAddRecFN.scala 121:16:chipyard.TestHarness.RocketConfig.fir@233577.4]
  assign _T_68 = doSubMags ? 53'h1fffffffffffff : 53'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@233579.4]
  assign _T_70 = {_T_66,_T_68}; // @[MulAddRecFN.scala 123:11:chipyard.TestHarness.RocketConfig.fir@233581.4]
  assign mainAlignedSigC = $signed(_T_70) >>> CAlignDist; // @[MulAddRecFN.scala 123:17:chipyard.TestHarness.RocketConfig.fir@233582.4]
  assign _T_71 = {rawC_sig, 2'h0}; // @[MulAddRecFN.scala 125:30:chipyard.TestHarness.RocketConfig.fir@233583.4]
  assign _T_74 = |_T_71[3:0]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233587.4]
  assign _T_76 = |_T_71[7:4]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233590.4]
  assign _T_78 = |_T_71[11:8]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233593.4]
  assign _T_80 = |_T_71[15:12]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233596.4]
  assign _T_82 = |_T_71[19:16]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233599.4]
  assign _T_84 = |_T_71[23:20]; // @[primitives.scala 121:54:chipyard.TestHarness.RocketConfig.fir@233602.4]
  assign _T_86 = |_T_71[26:24]; // @[primitives.scala 124:57:chipyard.TestHarness.RocketConfig.fir@233605.4]
  assign _T_92 = {_T_86,_T_84,_T_82,_T_80,_T_78,_T_76,_T_74}; // @[primitives.scala 125:20:chipyard.TestHarness.RocketConfig.fir@233612.4]
  assign _T_94 = -33'sh100000000 >>> CAlignDist[6:2]; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@233614.4]
  assign _T_110 = {_T_94[14],_T_94[15],_T_94[16],_T_94[17],_T_94[18],_T_94[19]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233630.4]
  assign _GEN_1 = {{1'd0}, _T_110}; // @[MulAddRecFN.scala 125:68:chipyard.TestHarness.RocketConfig.fir@233631.4]
  assign _T_111 = _T_92 & _GEN_1; // @[MulAddRecFN.scala 125:68:chipyard.TestHarness.RocketConfig.fir@233631.4]
  assign reduced4CExtra = |_T_111; // @[MulAddRecFN.scala 133:11:chipyard.TestHarness.RocketConfig.fir@233632.4]
  assign _T_114 = &mainAlignedSigC[2:0]; // @[MulAddRecFN.scala 137:39:chipyard.TestHarness.RocketConfig.fir@233635.4]
  assign _T_115 = ~reduced4CExtra; // @[MulAddRecFN.scala 137:47:chipyard.TestHarness.RocketConfig.fir@233636.4]
  assign _T_116 = _T_114 & _T_115; // @[MulAddRecFN.scala 137:44:chipyard.TestHarness.RocketConfig.fir@233637.4]
  assign _T_118 = |mainAlignedSigC[2:0]; // @[MulAddRecFN.scala 138:39:chipyard.TestHarness.RocketConfig.fir@233639.4]
  assign _T_119 = _T_118 | reduced4CExtra; // @[MulAddRecFN.scala 138:44:chipyard.TestHarness.RocketConfig.fir@233640.4]
  assign _T_120 = doSubMags ? _T_116 : _T_119; // @[MulAddRecFN.scala 136:16:chipyard.TestHarness.RocketConfig.fir@233641.4]
  assign _T_121 = mainAlignedSigC[77:3]; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233642.4]
  assign alignedSigC = {_T_121,_T_120}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@233643.4]
  assign _T_124 = ~rawA_sig[22]; // @[common.scala 81:49:chipyard.TestHarness.RocketConfig.fir@233649.4]
  assign _T_125 = rawA_isNaN & _T_124; // @[common.scala 81:46:chipyard.TestHarness.RocketConfig.fir@233650.4]
  assign _T_127 = ~rawB_sig[22]; // @[common.scala 81:49:chipyard.TestHarness.RocketConfig.fir@233652.4]
  assign _T_128 = rawB_isNaN & _T_127; // @[common.scala 81:46:chipyard.TestHarness.RocketConfig.fir@233653.4]
  assign _T_129 = _T_125 | _T_128; // @[MulAddRecFN.scala 149:32:chipyard.TestHarness.RocketConfig.fir@233654.4]
  assign _T_131 = ~rawC_sig[22]; // @[common.scala 81:49:chipyard.TestHarness.RocketConfig.fir@233656.4]
  assign _T_132 = rawC_isNaN & _T_131; // @[common.scala 81:46:chipyard.TestHarness.RocketConfig.fir@233657.4]
  assign _T_137 = $signed(sExpAlignedProd) - 11'sh18; // @[MulAddRecFN.scala 161:53:chipyard.TestHarness.RocketConfig.fir@233672.4]
  assign _T_138 = CIsDominant ? $signed({{1{rawC_sExp[9]}},rawC_sExp}) : $signed(_T_137); // @[MulAddRecFN.scala 161:12:chipyard.TestHarness.RocketConfig.fir@233673.4]
  assign io_mulAddA = rawA_sig[23:0]; // @[MulAddRecFN.scala 144:16:chipyard.TestHarness.RocketConfig.fir@233644.4]
  assign io_mulAddB = rawB_sig[23:0]; // @[MulAddRecFN.scala 145:16:chipyard.TestHarness.RocketConfig.fir@233645.4]
  assign io_mulAddC = alignedSigC[48:1]; // @[MulAddRecFN.scala 146:16:chipyard.TestHarness.RocketConfig.fir@233647.4]
  assign io_toPostMul_isSigNaNAny = _T_129 | _T_132; // @[MulAddRecFN.scala 148:30:chipyard.TestHarness.RocketConfig.fir@233659.4]
  assign io_toPostMul_isNaNAOrB = rawA_isNaN | rawB_isNaN; // @[MulAddRecFN.scala 151:28:chipyard.TestHarness.RocketConfig.fir@233661.4]
  assign io_toPostMul_isInfA = _T_4 & _T_8; // @[MulAddRecFN.scala 152:28:chipyard.TestHarness.RocketConfig.fir@233662.4]
  assign io_toPostMul_isZeroA = io_a[31:29] == 3'h0; // @[MulAddRecFN.scala 153:28:chipyard.TestHarness.RocketConfig.fir@233663.4]
  assign io_toPostMul_isInfB = _T_20 & _T_24; // @[MulAddRecFN.scala 154:28:chipyard.TestHarness.RocketConfig.fir@233664.4]
  assign io_toPostMul_isZeroB = io_b[31:29] == 3'h0; // @[MulAddRecFN.scala 155:28:chipyard.TestHarness.RocketConfig.fir@233665.4]
  assign io_toPostMul_signProd = _T_48 ^ io_op[1]; // @[MulAddRecFN.scala 156:28:chipyard.TestHarness.RocketConfig.fir@233666.4]
  assign io_toPostMul_isNaNC = _T_36 & io_c[29]; // @[MulAddRecFN.scala 157:28:chipyard.TestHarness.RocketConfig.fir@233667.4]
  assign io_toPostMul_isInfC = _T_36 & _T_40; // @[MulAddRecFN.scala 158:28:chipyard.TestHarness.RocketConfig.fir@233668.4]
  assign io_toPostMul_isZeroC = io_c[31:29] == 3'h0; // @[MulAddRecFN.scala 159:28:chipyard.TestHarness.RocketConfig.fir@233669.4]
  assign io_toPostMul_sExpSum = _T_138[9:0]; // @[MulAddRecFN.scala 160:28:chipyard.TestHarness.RocketConfig.fir@233674.4]
  assign io_toPostMul_doSubMags = _T_53 ^ io_op[0]; // @[MulAddRecFN.scala 162:28:chipyard.TestHarness.RocketConfig.fir@233675.4]
  assign io_toPostMul_CIsDominant = _T_44 & _T_61; // @[MulAddRecFN.scala 163:30:chipyard.TestHarness.RocketConfig.fir@233676.4]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[4:0]; // @[MulAddRecFN.scala 164:34:chipyard.TestHarness.RocketConfig.fir@233678.4]
  assign io_toPostMul_highAlignedSigC = alignedSigC[74:49]; // @[MulAddRecFN.scala 165:34:chipyard.TestHarness.RocketConfig.fir@233680.4]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:34:chipyard.TestHarness.RocketConfig.fir@233682.4]
endmodule
