module PMPChecker( // @[:chipyard.TestHarness.RocketConfig.fir@195823.2]
  input  [1:0]  io_prv, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_0_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [1:0]  io_pmp_0_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_0_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_0_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_0_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [29:0] io_pmp_0_addr, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [31:0] io_pmp_0_mask, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_1_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [1:0]  io_pmp_1_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_1_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_1_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_1_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [29:0] io_pmp_1_addr, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [31:0] io_pmp_1_mask, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_2_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [1:0]  io_pmp_2_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_2_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_2_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_2_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [29:0] io_pmp_2_addr, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [31:0] io_pmp_2_mask, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_3_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [1:0]  io_pmp_3_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_3_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_3_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_3_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [29:0] io_pmp_3_addr, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [31:0] io_pmp_3_mask, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_4_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [1:0]  io_pmp_4_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_4_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_4_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_4_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [29:0] io_pmp_4_addr, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [31:0] io_pmp_4_mask, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_5_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [1:0]  io_pmp_5_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_5_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_5_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_5_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [29:0] io_pmp_5_addr, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [31:0] io_pmp_5_mask, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_6_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [1:0]  io_pmp_6_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_6_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_6_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_6_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [29:0] io_pmp_6_addr, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [31:0] io_pmp_6_mask, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_7_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [1:0]  io_pmp_7_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_7_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_7_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input         io_pmp_7_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [29:0] io_pmp_7_addr, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [31:0] io_pmp_7_mask, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [31:0] io_addr, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  input  [1:0]  io_size, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  output        io_r, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  output        io_w, // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
  output        io_x // @[:chipyard.TestHarness.RocketConfig.fir@195826.4]
);
  wire  default_; // @[PMP.scala 157:56:chipyard.TestHarness.RocketConfig.fir@195828.4]
  wire [5:0] _T_3; // @[package.scala 189:77:chipyard.TestHarness.RocketConfig.fir@195852.4]
  wire [2:0] _T_5; // @[package.scala 189:46:chipyard.TestHarness.RocketConfig.fir@195854.4]
  wire [31:0] _GEN_0; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@195855.4]
  wire [31:0] _T_6; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@195855.4]
  wire [31:0] _T_8; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@195857.4]
  wire [31:0] _T_9; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@195858.4]
  wire [31:0] _T_10; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@195859.4]
  wire [31:0] _T_11; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@195860.4]
  wire [28:0] _T_14; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@195863.4]
  wire [28:0] _T_15; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@195864.4]
  wire [28:0] _T_16; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@195865.4]
  wire  _T_17; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@195866.4]
  wire [2:0] _T_25; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@195874.4]
  wire [2:0] _T_26; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@195875.4]
  wire [2:0] _T_27; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@195876.4]
  wire  _T_28; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@195877.4]
  wire  _T_29; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@195878.4]
  wire [31:0] _T_36; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@195885.4]
  wire [31:0] _T_37; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@195886.4]
  wire [31:0] _T_38; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@195887.4]
  wire [31:0] _T_39; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@195888.4]
  wire  _T_41; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@195890.4]
  wire [28:0] _T_48; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@195897.4]
  wire  _T_49; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@195898.4]
  wire [2:0] _T_51; // @[PMP.scala 84:42:chipyard.TestHarness.RocketConfig.fir@195900.4]
  wire  _T_57; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@195906.4]
  wire  _T_58; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@195907.4]
  wire  _T_59; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@195908.4]
  wire  _T_60; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@195909.4]
  wire  _T_67; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@195916.4]
  wire  _T_75; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@195924.4]
  wire  _T_83; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@195932.4]
  wire  _T_84; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@195933.4]
  wire  _T_85; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@195934.4]
  wire  _T_86; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@195935.4]
  wire  _T_87; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@195936.4]
  wire  _T_88; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@195937.4]
  wire  _T_89; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@195938.4]
  wire  _T_90; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@195939.4]
  wire [2:0] _T_109; // @[PMP.scala 125:125:chipyard.TestHarness.RocketConfig.fir@195958.4]
  wire [2:0] _T_110; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@195959.4]
  wire  _T_111; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@195960.4]
  wire  _T_112; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@195961.4]
  wire [2:0] _T_128; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@195977.4]
  wire  _T_129; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@195978.4]
  wire  _T_130; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@195979.4]
  wire  _T_131; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@195980.4]
  wire  _T_132; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@195981.4]
  wire [2:0] _T_134; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@195983.4]
  wire [2:0] _T_135; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@195984.4]
  wire  _T_136; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@195985.4]
  wire  _T_138; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@195987.4]
  wire  _T_190; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@196047.4]
  wire  _T_191; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@196048.4]
  wire  _T_192; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@196050.4]
  wire  _T_193; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@196051.4]
  wire  _T_194; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@196053.4]
  wire  _T_195; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@196054.4]
  wire  _T_196_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196056.4]
  wire  _T_196_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196056.4]
  wire  _T_196_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196056.4]
  wire [31:0] _T_202; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@196062.4]
  wire [28:0] _T_211; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196071.4]
  wire [28:0] _T_212; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196072.4]
  wire  _T_213; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196073.4]
  wire [2:0] _T_221; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@196081.4]
  wire [2:0] _T_222; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196082.4]
  wire [2:0] _T_223; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196083.4]
  wire  _T_224; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196084.4]
  wire  _T_225; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@196085.4]
  wire [31:0] _T_232; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@196092.4]
  wire [31:0] _T_233; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@196093.4]
  wire [31:0] _T_234; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@196094.4]
  wire [31:0] _T_235; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@196095.4]
  wire  _T_237; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@196097.4]
  wire [28:0] _T_244; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@196104.4]
  wire  _T_245; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@196105.4]
  wire  _T_253; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196113.4]
  wire  _T_254; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196114.4]
  wire  _T_255; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196115.4]
  wire  _T_256; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@196116.4]
  wire  _T_279; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196139.4]
  wire  _T_280; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196140.4]
  wire  _T_281; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196141.4]
  wire  _T_282; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@196142.4]
  wire  _T_283; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@196143.4]
  wire  _T_284; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@196144.4]
  wire  _T_285; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@196145.4]
  wire  _T_286; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@196146.4]
  wire [2:0] _T_306; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@196166.4]
  wire  _T_307; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@196167.4]
  wire  _T_308; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@196168.4]
  wire [2:0] _T_324; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@196184.4]
  wire  _T_325; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@196185.4]
  wire  _T_326; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@196186.4]
  wire  _T_327; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@196187.4]
  wire  _T_328; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@196188.4]
  wire [2:0] _T_330; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@196190.4]
  wire [2:0] _T_331; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@196191.4]
  wire  _T_332; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@196192.4]
  wire  _T_334; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@196194.4]
  wire  _T_386; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@196254.4]
  wire  _T_387; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@196255.4]
  wire  _T_388; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@196257.4]
  wire  _T_389; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@196258.4]
  wire  _T_390; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@196260.4]
  wire  _T_391; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@196261.4]
  wire  _T_392_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196263.4]
  wire  _T_392_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196263.4]
  wire  _T_392_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196263.4]
  wire [31:0] _T_398; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@196269.4]
  wire [28:0] _T_407; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196278.4]
  wire [28:0] _T_408; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196279.4]
  wire  _T_409; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196280.4]
  wire [2:0] _T_417; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@196288.4]
  wire [2:0] _T_418; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196289.4]
  wire [2:0] _T_419; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196290.4]
  wire  _T_420; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196291.4]
  wire  _T_421; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@196292.4]
  wire [31:0] _T_428; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@196299.4]
  wire [31:0] _T_429; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@196300.4]
  wire [31:0] _T_430; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@196301.4]
  wire [31:0] _T_431; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@196302.4]
  wire  _T_433; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@196304.4]
  wire [28:0] _T_440; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@196311.4]
  wire  _T_441; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@196312.4]
  wire  _T_449; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196320.4]
  wire  _T_450; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196321.4]
  wire  _T_451; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196322.4]
  wire  _T_452; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@196323.4]
  wire  _T_475; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196346.4]
  wire  _T_476; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196347.4]
  wire  _T_477; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196348.4]
  wire  _T_478; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@196349.4]
  wire  _T_479; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@196350.4]
  wire  _T_480; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@196351.4]
  wire  _T_481; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@196352.4]
  wire  _T_482; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@196353.4]
  wire [2:0] _T_502; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@196373.4]
  wire  _T_503; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@196374.4]
  wire  _T_504; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@196375.4]
  wire [2:0] _T_520; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@196391.4]
  wire  _T_521; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@196392.4]
  wire  _T_522; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@196393.4]
  wire  _T_523; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@196394.4]
  wire  _T_524; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@196395.4]
  wire [2:0] _T_526; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@196397.4]
  wire [2:0] _T_527; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@196398.4]
  wire  _T_528; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@196399.4]
  wire  _T_530; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@196401.4]
  wire  _T_582; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@196461.4]
  wire  _T_583; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@196462.4]
  wire  _T_584; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@196464.4]
  wire  _T_585; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@196465.4]
  wire  _T_586; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@196467.4]
  wire  _T_587; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@196468.4]
  wire  _T_588_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196470.4]
  wire  _T_588_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196470.4]
  wire  _T_588_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196470.4]
  wire [31:0] _T_594; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@196476.4]
  wire [28:0] _T_603; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196485.4]
  wire [28:0] _T_604; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196486.4]
  wire  _T_605; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196487.4]
  wire [2:0] _T_613; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@196495.4]
  wire [2:0] _T_614; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196496.4]
  wire [2:0] _T_615; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196497.4]
  wire  _T_616; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196498.4]
  wire  _T_617; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@196499.4]
  wire [31:0] _T_624; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@196506.4]
  wire [31:0] _T_625; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@196507.4]
  wire [31:0] _T_626; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@196508.4]
  wire [31:0] _T_627; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@196509.4]
  wire  _T_629; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@196511.4]
  wire [28:0] _T_636; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@196518.4]
  wire  _T_637; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@196519.4]
  wire  _T_645; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196527.4]
  wire  _T_646; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196528.4]
  wire  _T_647; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196529.4]
  wire  _T_648; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@196530.4]
  wire  _T_671; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196553.4]
  wire  _T_672; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196554.4]
  wire  _T_673; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196555.4]
  wire  _T_674; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@196556.4]
  wire  _T_675; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@196557.4]
  wire  _T_676; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@196558.4]
  wire  _T_677; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@196559.4]
  wire  _T_678; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@196560.4]
  wire [2:0] _T_698; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@196580.4]
  wire  _T_699; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@196581.4]
  wire  _T_700; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@196582.4]
  wire [2:0] _T_716; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@196598.4]
  wire  _T_717; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@196599.4]
  wire  _T_718; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@196600.4]
  wire  _T_719; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@196601.4]
  wire  _T_720; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@196602.4]
  wire [2:0] _T_722; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@196604.4]
  wire [2:0] _T_723; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@196605.4]
  wire  _T_724; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@196606.4]
  wire  _T_726; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@196608.4]
  wire  _T_778; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@196668.4]
  wire  _T_779; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@196669.4]
  wire  _T_780; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@196671.4]
  wire  _T_781; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@196672.4]
  wire  _T_782; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@196674.4]
  wire  _T_783; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@196675.4]
  wire  _T_784_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196677.4]
  wire  _T_784_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196677.4]
  wire  _T_784_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196677.4]
  wire [31:0] _T_790; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@196683.4]
  wire [28:0] _T_799; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196692.4]
  wire [28:0] _T_800; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196693.4]
  wire  _T_801; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196694.4]
  wire [2:0] _T_809; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@196702.4]
  wire [2:0] _T_810; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196703.4]
  wire [2:0] _T_811; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196704.4]
  wire  _T_812; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196705.4]
  wire  _T_813; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@196706.4]
  wire [31:0] _T_820; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@196713.4]
  wire [31:0] _T_821; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@196714.4]
  wire [31:0] _T_822; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@196715.4]
  wire [31:0] _T_823; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@196716.4]
  wire  _T_825; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@196718.4]
  wire [28:0] _T_832; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@196725.4]
  wire  _T_833; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@196726.4]
  wire  _T_841; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196734.4]
  wire  _T_842; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196735.4]
  wire  _T_843; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196736.4]
  wire  _T_844; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@196737.4]
  wire  _T_867; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196760.4]
  wire  _T_868; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196761.4]
  wire  _T_869; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196762.4]
  wire  _T_870; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@196763.4]
  wire  _T_871; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@196764.4]
  wire  _T_872; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@196765.4]
  wire  _T_873; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@196766.4]
  wire  _T_874; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@196767.4]
  wire [2:0] _T_894; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@196787.4]
  wire  _T_895; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@196788.4]
  wire  _T_896; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@196789.4]
  wire [2:0] _T_912; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@196805.4]
  wire  _T_913; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@196806.4]
  wire  _T_914; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@196807.4]
  wire  _T_915; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@196808.4]
  wire  _T_916; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@196809.4]
  wire [2:0] _T_918; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@196811.4]
  wire [2:0] _T_919; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@196812.4]
  wire  _T_920; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@196813.4]
  wire  _T_922; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@196815.4]
  wire  _T_974; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@196875.4]
  wire  _T_975; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@196876.4]
  wire  _T_976; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@196878.4]
  wire  _T_977; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@196879.4]
  wire  _T_978; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@196881.4]
  wire  _T_979; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@196882.4]
  wire  _T_980_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196884.4]
  wire  _T_980_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196884.4]
  wire  _T_980_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196884.4]
  wire [31:0] _T_986; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@196890.4]
  wire [28:0] _T_995; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196899.4]
  wire [28:0] _T_996; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196900.4]
  wire  _T_997; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196901.4]
  wire [2:0] _T_1005; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@196909.4]
  wire [2:0] _T_1006; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196910.4]
  wire [2:0] _T_1007; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196911.4]
  wire  _T_1008; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196912.4]
  wire  _T_1009; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@196913.4]
  wire [31:0] _T_1016; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@196920.4]
  wire [31:0] _T_1017; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@196921.4]
  wire [31:0] _T_1018; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@196922.4]
  wire [31:0] _T_1019; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@196923.4]
  wire  _T_1021; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@196925.4]
  wire [28:0] _T_1028; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@196932.4]
  wire  _T_1029; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@196933.4]
  wire  _T_1037; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196941.4]
  wire  _T_1038; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196942.4]
  wire  _T_1039; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196943.4]
  wire  _T_1040; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@196944.4]
  wire  _T_1063; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196967.4]
  wire  _T_1064; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196968.4]
  wire  _T_1065; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196969.4]
  wire  _T_1066; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@196970.4]
  wire  _T_1067; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@196971.4]
  wire  _T_1068; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@196972.4]
  wire  _T_1069; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@196973.4]
  wire  _T_1070; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@196974.4]
  wire [2:0] _T_1090; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@196994.4]
  wire  _T_1091; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@196995.4]
  wire  _T_1092; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@196996.4]
  wire [2:0] _T_1108; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@197012.4]
  wire  _T_1109; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@197013.4]
  wire  _T_1110; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@197014.4]
  wire  _T_1111; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@197015.4]
  wire  _T_1112; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@197016.4]
  wire [2:0] _T_1114; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@197018.4]
  wire [2:0] _T_1115; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@197019.4]
  wire  _T_1116; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@197020.4]
  wire  _T_1118; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@197022.4]
  wire  _T_1170; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@197082.4]
  wire  _T_1171; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@197083.4]
  wire  _T_1172; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@197085.4]
  wire  _T_1173; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@197086.4]
  wire  _T_1174; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@197088.4]
  wire  _T_1175; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@197089.4]
  wire  _T_1176_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@197091.4]
  wire  _T_1176_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@197091.4]
  wire  _T_1176_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@197091.4]
  wire [31:0] _T_1182; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@197097.4]
  wire [28:0] _T_1191; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@197106.4]
  wire [28:0] _T_1192; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@197107.4]
  wire  _T_1193; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@197108.4]
  wire [2:0] _T_1201; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@197116.4]
  wire [2:0] _T_1202; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@197117.4]
  wire [2:0] _T_1203; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@197118.4]
  wire  _T_1204; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@197119.4]
  wire  _T_1205; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@197120.4]
  wire [31:0] _T_1212; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@197127.4]
  wire [31:0] _T_1213; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@197128.4]
  wire [31:0] _T_1214; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@197129.4]
  wire [31:0] _T_1215; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@197130.4]
  wire  _T_1217; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@197132.4]
  wire [28:0] _T_1224; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@197139.4]
  wire  _T_1225; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@197140.4]
  wire  _T_1233; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@197148.4]
  wire  _T_1234; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@197149.4]
  wire  _T_1235; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@197150.4]
  wire  _T_1236; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@197151.4]
  wire  _T_1259; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@197174.4]
  wire  _T_1260; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@197175.4]
  wire  _T_1261; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@197176.4]
  wire  _T_1262; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@197177.4]
  wire  _T_1263; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@197178.4]
  wire  _T_1264; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@197179.4]
  wire  _T_1265; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@197180.4]
  wire  _T_1266; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@197181.4]
  wire [2:0] _T_1286; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@197201.4]
  wire  _T_1287; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@197202.4]
  wire  _T_1288; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@197203.4]
  wire [2:0] _T_1304; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@197219.4]
  wire  _T_1305; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@197220.4]
  wire  _T_1306; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@197221.4]
  wire  _T_1307; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@197222.4]
  wire  _T_1308; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@197223.4]
  wire [2:0] _T_1310; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@197225.4]
  wire [2:0] _T_1311; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@197226.4]
  wire  _T_1312; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@197227.4]
  wire  _T_1314; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@197229.4]
  wire  _T_1366; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@197289.4]
  wire  _T_1367; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@197290.4]
  wire  _T_1368; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@197292.4]
  wire  _T_1369; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@197293.4]
  wire  _T_1370; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@197295.4]
  wire  _T_1371; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@197296.4]
  wire  _T_1372_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@197298.4]
  wire  _T_1372_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@197298.4]
  wire  _T_1372_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@197298.4]
  wire [31:0] _T_1378; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@197304.4]
  wire [28:0] _T_1387; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@197313.4]
  wire [28:0] _T_1388; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@197314.4]
  wire  _T_1389; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@197315.4]
  wire [2:0] _T_1397; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@197323.4]
  wire [2:0] _T_1398; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@197324.4]
  wire [2:0] _T_1399; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@197325.4]
  wire  _T_1400; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@197326.4]
  wire  _T_1401; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@197327.4]
  wire  _T_1455; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@197381.4]
  wire  _T_1456; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@197382.4]
  wire  _T_1457; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@197383.4]
  wire  _T_1459; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@197385.4]
  wire  _T_1460; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@197386.4]
  wire  _T_1461; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@197387.4]
  wire  _T_1462; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@197388.4]
  wire [2:0] _T_1500; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@197426.4]
  wire  _T_1501; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@197427.4]
  wire  _T_1502; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@197428.4]
  wire  _T_1504; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@197430.4]
  wire [2:0] _T_1506; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@197432.4]
  wire [2:0] _T_1507; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@197433.4]
  wire  _T_1508; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@197434.4]
  wire  _T_1510; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@197436.4]
  wire  _T_1562; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@197496.4]
  wire  _T_1563; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@197497.4]
  wire  _T_1564; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@197499.4]
  wire  _T_1565; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@197500.4]
  wire  _T_1566; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@197502.4]
  wire  _T_1567; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@197503.4]
  assign default_ = io_prv > 2'h1; // @[PMP.scala 157:56:chipyard.TestHarness.RocketConfig.fir@195828.4]
  assign _T_3 = 6'h7 << io_size; // @[package.scala 189:77:chipyard.TestHarness.RocketConfig.fir@195852.4]
  assign _T_5 = ~_T_3[2:0]; // @[package.scala 189:46:chipyard.TestHarness.RocketConfig.fir@195854.4]
  assign _GEN_0 = {{29'd0}, _T_5}; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@195855.4]
  assign _T_6 = io_pmp_7_mask | _GEN_0; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@195855.4]
  assign _T_8 = {io_pmp_7_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@195857.4]
  assign _T_9 = ~_T_8; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@195858.4]
  assign _T_10 = _T_9 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@195859.4]
  assign _T_11 = ~_T_10; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@195860.4]
  assign _T_14 = io_addr[31:3] ^ _T_11[31:3]; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@195863.4]
  assign _T_15 = ~io_pmp_7_mask[31:3]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@195864.4]
  assign _T_16 = _T_14 & _T_15; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@195865.4]
  assign _T_17 = _T_16 == 29'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@195866.4]
  assign _T_25 = io_addr[2:0] ^ _T_11[2:0]; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@195874.4]
  assign _T_26 = ~_T_6[2:0]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@195875.4]
  assign _T_27 = _T_25 & _T_26; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@195876.4]
  assign _T_28 = _T_27 == 3'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@195877.4]
  assign _T_29 = _T_17 & _T_28; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@195878.4]
  assign _T_36 = {io_pmp_6_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@195885.4]
  assign _T_37 = ~_T_36; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@195886.4]
  assign _T_38 = _T_37 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@195887.4]
  assign _T_39 = ~_T_38; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@195888.4]
  assign _T_41 = io_addr[31:3] < _T_39[31:3]; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@195890.4]
  assign _T_48 = io_addr[31:3] ^ _T_39[31:3]; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@195897.4]
  assign _T_49 = _T_48 == 29'h0; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@195898.4]
  assign _T_51 = io_addr[2:0] | _T_5; // @[PMP.scala 84:42:chipyard.TestHarness.RocketConfig.fir@195900.4]
  assign _T_57 = _T_51 < _T_39[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@195906.4]
  assign _T_58 = _T_49 & _T_57; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@195907.4]
  assign _T_59 = _T_41 | _T_58; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@195908.4]
  assign _T_60 = ~_T_59; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@195909.4]
  assign _T_67 = io_addr[31:3] < _T_11[31:3]; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@195916.4]
  assign _T_75 = _T_14 == 29'h0; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@195924.4]
  assign _T_83 = io_addr[2:0] < _T_11[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@195932.4]
  assign _T_84 = _T_75 & _T_83; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@195933.4]
  assign _T_85 = _T_67 | _T_84; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@195934.4]
  assign _T_86 = _T_60 & _T_85; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@195935.4]
  assign _T_87 = io_pmp_7_cfg_a[0] & _T_86; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@195936.4]
  assign _T_88 = io_pmp_7_cfg_a[1] ? _T_29 : _T_87; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@195937.4]
  assign _T_89 = ~io_pmp_7_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@195938.4]
  assign _T_90 = default_ & _T_89; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@195939.4]
  assign _T_109 = ~io_addr[2:0]; // @[PMP.scala 125:125:chipyard.TestHarness.RocketConfig.fir@195958.4]
  assign _T_110 = _T_39[2:0] & _T_109; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@195959.4]
  assign _T_111 = _T_110 != 3'h0; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@195960.4]
  assign _T_112 = _T_49 & _T_111; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@195961.4]
  assign _T_128 = _T_11[2:0] & _T_51; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@195977.4]
  assign _T_129 = _T_128 != 3'h0; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@195978.4]
  assign _T_130 = _T_75 & _T_129; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@195979.4]
  assign _T_131 = _T_112 | _T_130; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@195980.4]
  assign _T_132 = ~_T_131; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@195981.4]
  assign _T_134 = ~io_pmp_7_mask[2:0]; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@195983.4]
  assign _T_135 = _T_5 & _T_134; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@195984.4]
  assign _T_136 = _T_135 == 3'h0; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@195985.4]
  assign _T_138 = io_pmp_7_cfg_a[1] ? _T_136 : _T_132; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@195987.4]
  assign _T_190 = io_pmp_7_cfg_r | _T_90; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@196047.4]
  assign _T_191 = _T_138 & _T_190; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@196048.4]
  assign _T_192 = io_pmp_7_cfg_w | _T_90; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@196050.4]
  assign _T_193 = _T_138 & _T_192; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@196051.4]
  assign _T_194 = io_pmp_7_cfg_x | _T_90; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@196053.4]
  assign _T_195 = _T_138 & _T_194; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@196054.4]
  assign _T_196_cfg_x = _T_88 ? _T_195 : default_; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196056.4]
  assign _T_196_cfg_w = _T_88 ? _T_193 : default_; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196056.4]
  assign _T_196_cfg_r = _T_88 ? _T_191 : default_; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196056.4]
  assign _T_202 = io_pmp_6_mask | _GEN_0; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@196062.4]
  assign _T_211 = ~io_pmp_6_mask[31:3]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196071.4]
  assign _T_212 = _T_48 & _T_211; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196072.4]
  assign _T_213 = _T_212 == 29'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196073.4]
  assign _T_221 = io_addr[2:0] ^ _T_39[2:0]; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@196081.4]
  assign _T_222 = ~_T_202[2:0]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196082.4]
  assign _T_223 = _T_221 & _T_222; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196083.4]
  assign _T_224 = _T_223 == 3'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196084.4]
  assign _T_225 = _T_213 & _T_224; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@196085.4]
  assign _T_232 = {io_pmp_5_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@196092.4]
  assign _T_233 = ~_T_232; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@196093.4]
  assign _T_234 = _T_233 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@196094.4]
  assign _T_235 = ~_T_234; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@196095.4]
  assign _T_237 = io_addr[31:3] < _T_235[31:3]; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@196097.4]
  assign _T_244 = io_addr[31:3] ^ _T_235[31:3]; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@196104.4]
  assign _T_245 = _T_244 == 29'h0; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@196105.4]
  assign _T_253 = _T_51 < _T_235[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196113.4]
  assign _T_254 = _T_245 & _T_253; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196114.4]
  assign _T_255 = _T_237 | _T_254; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196115.4]
  assign _T_256 = ~_T_255; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@196116.4]
  assign _T_279 = io_addr[2:0] < _T_39[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196139.4]
  assign _T_280 = _T_49 & _T_279; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196140.4]
  assign _T_281 = _T_41 | _T_280; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196141.4]
  assign _T_282 = _T_256 & _T_281; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@196142.4]
  assign _T_283 = io_pmp_6_cfg_a[0] & _T_282; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@196143.4]
  assign _T_284 = io_pmp_6_cfg_a[1] ? _T_225 : _T_283; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@196144.4]
  assign _T_285 = ~io_pmp_6_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@196145.4]
  assign _T_286 = default_ & _T_285; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@196146.4]
  assign _T_306 = _T_235[2:0] & _T_109; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@196166.4]
  assign _T_307 = _T_306 != 3'h0; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@196167.4]
  assign _T_308 = _T_245 & _T_307; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@196168.4]
  assign _T_324 = _T_39[2:0] & _T_51; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@196184.4]
  assign _T_325 = _T_324 != 3'h0; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@196185.4]
  assign _T_326 = _T_49 & _T_325; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@196186.4]
  assign _T_327 = _T_308 | _T_326; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@196187.4]
  assign _T_328 = ~_T_327; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@196188.4]
  assign _T_330 = ~io_pmp_6_mask[2:0]; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@196190.4]
  assign _T_331 = _T_5 & _T_330; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@196191.4]
  assign _T_332 = _T_331 == 3'h0; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@196192.4]
  assign _T_334 = io_pmp_6_cfg_a[1] ? _T_332 : _T_328; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@196194.4]
  assign _T_386 = io_pmp_6_cfg_r | _T_286; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@196254.4]
  assign _T_387 = _T_334 & _T_386; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@196255.4]
  assign _T_388 = io_pmp_6_cfg_w | _T_286; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@196257.4]
  assign _T_389 = _T_334 & _T_388; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@196258.4]
  assign _T_390 = io_pmp_6_cfg_x | _T_286; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@196260.4]
  assign _T_391 = _T_334 & _T_390; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@196261.4]
  assign _T_392_cfg_x = _T_284 ? _T_391 : _T_196_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196263.4]
  assign _T_392_cfg_w = _T_284 ? _T_389 : _T_196_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196263.4]
  assign _T_392_cfg_r = _T_284 ? _T_387 : _T_196_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196263.4]
  assign _T_398 = io_pmp_5_mask | _GEN_0; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@196269.4]
  assign _T_407 = ~io_pmp_5_mask[31:3]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196278.4]
  assign _T_408 = _T_244 & _T_407; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196279.4]
  assign _T_409 = _T_408 == 29'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196280.4]
  assign _T_417 = io_addr[2:0] ^ _T_235[2:0]; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@196288.4]
  assign _T_418 = ~_T_398[2:0]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196289.4]
  assign _T_419 = _T_417 & _T_418; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196290.4]
  assign _T_420 = _T_419 == 3'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196291.4]
  assign _T_421 = _T_409 & _T_420; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@196292.4]
  assign _T_428 = {io_pmp_4_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@196299.4]
  assign _T_429 = ~_T_428; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@196300.4]
  assign _T_430 = _T_429 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@196301.4]
  assign _T_431 = ~_T_430; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@196302.4]
  assign _T_433 = io_addr[31:3] < _T_431[31:3]; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@196304.4]
  assign _T_440 = io_addr[31:3] ^ _T_431[31:3]; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@196311.4]
  assign _T_441 = _T_440 == 29'h0; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@196312.4]
  assign _T_449 = _T_51 < _T_431[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196320.4]
  assign _T_450 = _T_441 & _T_449; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196321.4]
  assign _T_451 = _T_433 | _T_450; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196322.4]
  assign _T_452 = ~_T_451; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@196323.4]
  assign _T_475 = io_addr[2:0] < _T_235[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196346.4]
  assign _T_476 = _T_245 & _T_475; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196347.4]
  assign _T_477 = _T_237 | _T_476; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196348.4]
  assign _T_478 = _T_452 & _T_477; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@196349.4]
  assign _T_479 = io_pmp_5_cfg_a[0] & _T_478; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@196350.4]
  assign _T_480 = io_pmp_5_cfg_a[1] ? _T_421 : _T_479; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@196351.4]
  assign _T_481 = ~io_pmp_5_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@196352.4]
  assign _T_482 = default_ & _T_481; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@196353.4]
  assign _T_502 = _T_431[2:0] & _T_109; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@196373.4]
  assign _T_503 = _T_502 != 3'h0; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@196374.4]
  assign _T_504 = _T_441 & _T_503; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@196375.4]
  assign _T_520 = _T_235[2:0] & _T_51; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@196391.4]
  assign _T_521 = _T_520 != 3'h0; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@196392.4]
  assign _T_522 = _T_245 & _T_521; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@196393.4]
  assign _T_523 = _T_504 | _T_522; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@196394.4]
  assign _T_524 = ~_T_523; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@196395.4]
  assign _T_526 = ~io_pmp_5_mask[2:0]; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@196397.4]
  assign _T_527 = _T_5 & _T_526; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@196398.4]
  assign _T_528 = _T_527 == 3'h0; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@196399.4]
  assign _T_530 = io_pmp_5_cfg_a[1] ? _T_528 : _T_524; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@196401.4]
  assign _T_582 = io_pmp_5_cfg_r | _T_482; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@196461.4]
  assign _T_583 = _T_530 & _T_582; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@196462.4]
  assign _T_584 = io_pmp_5_cfg_w | _T_482; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@196464.4]
  assign _T_585 = _T_530 & _T_584; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@196465.4]
  assign _T_586 = io_pmp_5_cfg_x | _T_482; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@196467.4]
  assign _T_587 = _T_530 & _T_586; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@196468.4]
  assign _T_588_cfg_x = _T_480 ? _T_587 : _T_392_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196470.4]
  assign _T_588_cfg_w = _T_480 ? _T_585 : _T_392_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196470.4]
  assign _T_588_cfg_r = _T_480 ? _T_583 : _T_392_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196470.4]
  assign _T_594 = io_pmp_4_mask | _GEN_0; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@196476.4]
  assign _T_603 = ~io_pmp_4_mask[31:3]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196485.4]
  assign _T_604 = _T_440 & _T_603; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196486.4]
  assign _T_605 = _T_604 == 29'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196487.4]
  assign _T_613 = io_addr[2:0] ^ _T_431[2:0]; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@196495.4]
  assign _T_614 = ~_T_594[2:0]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196496.4]
  assign _T_615 = _T_613 & _T_614; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196497.4]
  assign _T_616 = _T_615 == 3'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196498.4]
  assign _T_617 = _T_605 & _T_616; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@196499.4]
  assign _T_624 = {io_pmp_3_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@196506.4]
  assign _T_625 = ~_T_624; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@196507.4]
  assign _T_626 = _T_625 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@196508.4]
  assign _T_627 = ~_T_626; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@196509.4]
  assign _T_629 = io_addr[31:3] < _T_627[31:3]; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@196511.4]
  assign _T_636 = io_addr[31:3] ^ _T_627[31:3]; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@196518.4]
  assign _T_637 = _T_636 == 29'h0; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@196519.4]
  assign _T_645 = _T_51 < _T_627[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196527.4]
  assign _T_646 = _T_637 & _T_645; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196528.4]
  assign _T_647 = _T_629 | _T_646; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196529.4]
  assign _T_648 = ~_T_647; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@196530.4]
  assign _T_671 = io_addr[2:0] < _T_431[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196553.4]
  assign _T_672 = _T_441 & _T_671; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196554.4]
  assign _T_673 = _T_433 | _T_672; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196555.4]
  assign _T_674 = _T_648 & _T_673; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@196556.4]
  assign _T_675 = io_pmp_4_cfg_a[0] & _T_674; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@196557.4]
  assign _T_676 = io_pmp_4_cfg_a[1] ? _T_617 : _T_675; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@196558.4]
  assign _T_677 = ~io_pmp_4_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@196559.4]
  assign _T_678 = default_ & _T_677; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@196560.4]
  assign _T_698 = _T_627[2:0] & _T_109; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@196580.4]
  assign _T_699 = _T_698 != 3'h0; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@196581.4]
  assign _T_700 = _T_637 & _T_699; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@196582.4]
  assign _T_716 = _T_431[2:0] & _T_51; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@196598.4]
  assign _T_717 = _T_716 != 3'h0; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@196599.4]
  assign _T_718 = _T_441 & _T_717; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@196600.4]
  assign _T_719 = _T_700 | _T_718; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@196601.4]
  assign _T_720 = ~_T_719; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@196602.4]
  assign _T_722 = ~io_pmp_4_mask[2:0]; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@196604.4]
  assign _T_723 = _T_5 & _T_722; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@196605.4]
  assign _T_724 = _T_723 == 3'h0; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@196606.4]
  assign _T_726 = io_pmp_4_cfg_a[1] ? _T_724 : _T_720; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@196608.4]
  assign _T_778 = io_pmp_4_cfg_r | _T_678; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@196668.4]
  assign _T_779 = _T_726 & _T_778; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@196669.4]
  assign _T_780 = io_pmp_4_cfg_w | _T_678; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@196671.4]
  assign _T_781 = _T_726 & _T_780; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@196672.4]
  assign _T_782 = io_pmp_4_cfg_x | _T_678; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@196674.4]
  assign _T_783 = _T_726 & _T_782; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@196675.4]
  assign _T_784_cfg_x = _T_676 ? _T_783 : _T_588_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196677.4]
  assign _T_784_cfg_w = _T_676 ? _T_781 : _T_588_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196677.4]
  assign _T_784_cfg_r = _T_676 ? _T_779 : _T_588_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196677.4]
  assign _T_790 = io_pmp_3_mask | _GEN_0; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@196683.4]
  assign _T_799 = ~io_pmp_3_mask[31:3]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196692.4]
  assign _T_800 = _T_636 & _T_799; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196693.4]
  assign _T_801 = _T_800 == 29'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196694.4]
  assign _T_809 = io_addr[2:0] ^ _T_627[2:0]; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@196702.4]
  assign _T_810 = ~_T_790[2:0]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196703.4]
  assign _T_811 = _T_809 & _T_810; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196704.4]
  assign _T_812 = _T_811 == 3'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196705.4]
  assign _T_813 = _T_801 & _T_812; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@196706.4]
  assign _T_820 = {io_pmp_2_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@196713.4]
  assign _T_821 = ~_T_820; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@196714.4]
  assign _T_822 = _T_821 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@196715.4]
  assign _T_823 = ~_T_822; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@196716.4]
  assign _T_825 = io_addr[31:3] < _T_823[31:3]; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@196718.4]
  assign _T_832 = io_addr[31:3] ^ _T_823[31:3]; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@196725.4]
  assign _T_833 = _T_832 == 29'h0; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@196726.4]
  assign _T_841 = _T_51 < _T_823[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196734.4]
  assign _T_842 = _T_833 & _T_841; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196735.4]
  assign _T_843 = _T_825 | _T_842; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196736.4]
  assign _T_844 = ~_T_843; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@196737.4]
  assign _T_867 = io_addr[2:0] < _T_627[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196760.4]
  assign _T_868 = _T_637 & _T_867; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196761.4]
  assign _T_869 = _T_629 | _T_868; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196762.4]
  assign _T_870 = _T_844 & _T_869; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@196763.4]
  assign _T_871 = io_pmp_3_cfg_a[0] & _T_870; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@196764.4]
  assign _T_872 = io_pmp_3_cfg_a[1] ? _T_813 : _T_871; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@196765.4]
  assign _T_873 = ~io_pmp_3_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@196766.4]
  assign _T_874 = default_ & _T_873; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@196767.4]
  assign _T_894 = _T_823[2:0] & _T_109; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@196787.4]
  assign _T_895 = _T_894 != 3'h0; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@196788.4]
  assign _T_896 = _T_833 & _T_895; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@196789.4]
  assign _T_912 = _T_627[2:0] & _T_51; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@196805.4]
  assign _T_913 = _T_912 != 3'h0; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@196806.4]
  assign _T_914 = _T_637 & _T_913; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@196807.4]
  assign _T_915 = _T_896 | _T_914; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@196808.4]
  assign _T_916 = ~_T_915; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@196809.4]
  assign _T_918 = ~io_pmp_3_mask[2:0]; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@196811.4]
  assign _T_919 = _T_5 & _T_918; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@196812.4]
  assign _T_920 = _T_919 == 3'h0; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@196813.4]
  assign _T_922 = io_pmp_3_cfg_a[1] ? _T_920 : _T_916; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@196815.4]
  assign _T_974 = io_pmp_3_cfg_r | _T_874; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@196875.4]
  assign _T_975 = _T_922 & _T_974; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@196876.4]
  assign _T_976 = io_pmp_3_cfg_w | _T_874; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@196878.4]
  assign _T_977 = _T_922 & _T_976; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@196879.4]
  assign _T_978 = io_pmp_3_cfg_x | _T_874; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@196881.4]
  assign _T_979 = _T_922 & _T_978; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@196882.4]
  assign _T_980_cfg_x = _T_872 ? _T_979 : _T_784_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196884.4]
  assign _T_980_cfg_w = _T_872 ? _T_977 : _T_784_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196884.4]
  assign _T_980_cfg_r = _T_872 ? _T_975 : _T_784_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@196884.4]
  assign _T_986 = io_pmp_2_mask | _GEN_0; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@196890.4]
  assign _T_995 = ~io_pmp_2_mask[31:3]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196899.4]
  assign _T_996 = _T_832 & _T_995; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196900.4]
  assign _T_997 = _T_996 == 29'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196901.4]
  assign _T_1005 = io_addr[2:0] ^ _T_823[2:0]; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@196909.4]
  assign _T_1006 = ~_T_986[2:0]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@196910.4]
  assign _T_1007 = _T_1005 & _T_1006; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@196911.4]
  assign _T_1008 = _T_1007 == 3'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@196912.4]
  assign _T_1009 = _T_997 & _T_1008; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@196913.4]
  assign _T_1016 = {io_pmp_1_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@196920.4]
  assign _T_1017 = ~_T_1016; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@196921.4]
  assign _T_1018 = _T_1017 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@196922.4]
  assign _T_1019 = ~_T_1018; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@196923.4]
  assign _T_1021 = io_addr[31:3] < _T_1019[31:3]; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@196925.4]
  assign _T_1028 = io_addr[31:3] ^ _T_1019[31:3]; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@196932.4]
  assign _T_1029 = _T_1028 == 29'h0; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@196933.4]
  assign _T_1037 = _T_51 < _T_1019[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196941.4]
  assign _T_1038 = _T_1029 & _T_1037; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196942.4]
  assign _T_1039 = _T_1021 | _T_1038; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196943.4]
  assign _T_1040 = ~_T_1039; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@196944.4]
  assign _T_1063 = io_addr[2:0] < _T_823[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@196967.4]
  assign _T_1064 = _T_833 & _T_1063; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@196968.4]
  assign _T_1065 = _T_825 | _T_1064; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@196969.4]
  assign _T_1066 = _T_1040 & _T_1065; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@196970.4]
  assign _T_1067 = io_pmp_2_cfg_a[0] & _T_1066; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@196971.4]
  assign _T_1068 = io_pmp_2_cfg_a[1] ? _T_1009 : _T_1067; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@196972.4]
  assign _T_1069 = ~io_pmp_2_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@196973.4]
  assign _T_1070 = default_ & _T_1069; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@196974.4]
  assign _T_1090 = _T_1019[2:0] & _T_109; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@196994.4]
  assign _T_1091 = _T_1090 != 3'h0; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@196995.4]
  assign _T_1092 = _T_1029 & _T_1091; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@196996.4]
  assign _T_1108 = _T_823[2:0] & _T_51; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@197012.4]
  assign _T_1109 = _T_1108 != 3'h0; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@197013.4]
  assign _T_1110 = _T_833 & _T_1109; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@197014.4]
  assign _T_1111 = _T_1092 | _T_1110; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@197015.4]
  assign _T_1112 = ~_T_1111; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@197016.4]
  assign _T_1114 = ~io_pmp_2_mask[2:0]; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@197018.4]
  assign _T_1115 = _T_5 & _T_1114; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@197019.4]
  assign _T_1116 = _T_1115 == 3'h0; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@197020.4]
  assign _T_1118 = io_pmp_2_cfg_a[1] ? _T_1116 : _T_1112; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@197022.4]
  assign _T_1170 = io_pmp_2_cfg_r | _T_1070; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@197082.4]
  assign _T_1171 = _T_1118 & _T_1170; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@197083.4]
  assign _T_1172 = io_pmp_2_cfg_w | _T_1070; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@197085.4]
  assign _T_1173 = _T_1118 & _T_1172; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@197086.4]
  assign _T_1174 = io_pmp_2_cfg_x | _T_1070; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@197088.4]
  assign _T_1175 = _T_1118 & _T_1174; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@197089.4]
  assign _T_1176_cfg_x = _T_1068 ? _T_1175 : _T_980_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@197091.4]
  assign _T_1176_cfg_w = _T_1068 ? _T_1173 : _T_980_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@197091.4]
  assign _T_1176_cfg_r = _T_1068 ? _T_1171 : _T_980_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@197091.4]
  assign _T_1182 = io_pmp_1_mask | _GEN_0; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@197097.4]
  assign _T_1191 = ~io_pmp_1_mask[31:3]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@197106.4]
  assign _T_1192 = _T_1028 & _T_1191; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@197107.4]
  assign _T_1193 = _T_1192 == 29'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@197108.4]
  assign _T_1201 = io_addr[2:0] ^ _T_1019[2:0]; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@197116.4]
  assign _T_1202 = ~_T_1182[2:0]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@197117.4]
  assign _T_1203 = _T_1201 & _T_1202; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@197118.4]
  assign _T_1204 = _T_1203 == 3'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@197119.4]
  assign _T_1205 = _T_1193 & _T_1204; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@197120.4]
  assign _T_1212 = {io_pmp_0_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@197127.4]
  assign _T_1213 = ~_T_1212; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@197128.4]
  assign _T_1214 = _T_1213 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@197129.4]
  assign _T_1215 = ~_T_1214; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@197130.4]
  assign _T_1217 = io_addr[31:3] < _T_1215[31:3]; // @[PMP.scala 82:39:chipyard.TestHarness.RocketConfig.fir@197132.4]
  assign _T_1224 = io_addr[31:3] ^ _T_1215[31:3]; // @[PMP.scala 83:41:chipyard.TestHarness.RocketConfig.fir@197139.4]
  assign _T_1225 = _T_1224 == 29'h0; // @[PMP.scala 83:69:chipyard.TestHarness.RocketConfig.fir@197140.4]
  assign _T_1233 = _T_51 < _T_1215[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@197148.4]
  assign _T_1234 = _T_1225 & _T_1233; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@197149.4]
  assign _T_1235 = _T_1217 | _T_1234; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@197150.4]
  assign _T_1236 = ~_T_1235; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@197151.4]
  assign _T_1259 = io_addr[2:0] < _T_1019[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@197174.4]
  assign _T_1260 = _T_1029 & _T_1259; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@197175.4]
  assign _T_1261 = _T_1021 | _T_1260; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@197176.4]
  assign _T_1262 = _T_1236 & _T_1261; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@197177.4]
  assign _T_1263 = io_pmp_1_cfg_a[0] & _T_1262; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@197178.4]
  assign _T_1264 = io_pmp_1_cfg_a[1] ? _T_1205 : _T_1263; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@197179.4]
  assign _T_1265 = ~io_pmp_1_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@197180.4]
  assign _T_1266 = default_ & _T_1265; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@197181.4]
  assign _T_1286 = _T_1215[2:0] & _T_109; // @[PMP.scala 125:123:chipyard.TestHarness.RocketConfig.fir@197201.4]
  assign _T_1287 = _T_1286 != 3'h0; // @[PMP.scala 125:145:chipyard.TestHarness.RocketConfig.fir@197202.4]
  assign _T_1288 = _T_1225 & _T_1287; // @[PMP.scala 125:88:chipyard.TestHarness.RocketConfig.fir@197203.4]
  assign _T_1304 = _T_1019[2:0] & _T_51; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@197219.4]
  assign _T_1305 = _T_1304 != 3'h0; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@197220.4]
  assign _T_1306 = _T_1029 & _T_1305; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@197221.4]
  assign _T_1307 = _T_1288 | _T_1306; // @[PMP.scala 127:46:chipyard.TestHarness.RocketConfig.fir@197222.4]
  assign _T_1308 = ~_T_1307; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@197223.4]
  assign _T_1310 = ~io_pmp_1_mask[2:0]; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@197225.4]
  assign _T_1311 = _T_5 & _T_1310; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@197226.4]
  assign _T_1312 = _T_1311 == 3'h0; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@197227.4]
  assign _T_1314 = io_pmp_1_cfg_a[1] ? _T_1312 : _T_1308; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@197229.4]
  assign _T_1366 = io_pmp_1_cfg_r | _T_1266; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@197289.4]
  assign _T_1367 = _T_1314 & _T_1366; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@197290.4]
  assign _T_1368 = io_pmp_1_cfg_w | _T_1266; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@197292.4]
  assign _T_1369 = _T_1314 & _T_1368; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@197293.4]
  assign _T_1370 = io_pmp_1_cfg_x | _T_1266; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@197295.4]
  assign _T_1371 = _T_1314 & _T_1370; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@197296.4]
  assign _T_1372_cfg_x = _T_1264 ? _T_1371 : _T_1176_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@197298.4]
  assign _T_1372_cfg_w = _T_1264 ? _T_1369 : _T_1176_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@197298.4]
  assign _T_1372_cfg_r = _T_1264 ? _T_1367 : _T_1176_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@197298.4]
  assign _T_1378 = io_pmp_0_mask | _GEN_0; // @[PMP.scala 70:26:chipyard.TestHarness.RocketConfig.fir@197304.4]
  assign _T_1387 = ~io_pmp_0_mask[31:3]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@197313.4]
  assign _T_1388 = _T_1224 & _T_1387; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@197314.4]
  assign _T_1389 = _T_1388 == 29'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@197315.4]
  assign _T_1397 = io_addr[2:0] ^ _T_1215[2:0]; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@197323.4]
  assign _T_1398 = ~_T_1378[2:0]; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@197324.4]
  assign _T_1399 = _T_1397 & _T_1398; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@197325.4]
  assign _T_1400 = _T_1399 == 3'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@197326.4]
  assign _T_1401 = _T_1389 & _T_1400; // @[PMP.scala 73:16:chipyard.TestHarness.RocketConfig.fir@197327.4]
  assign _T_1455 = io_addr[2:0] < _T_1215[2:0]; // @[PMP.scala 84:53:chipyard.TestHarness.RocketConfig.fir@197381.4]
  assign _T_1456 = _T_1225 & _T_1455; // @[PMP.scala 85:30:chipyard.TestHarness.RocketConfig.fir@197382.4]
  assign _T_1457 = _T_1217 | _T_1456; // @[PMP.scala 85:16:chipyard.TestHarness.RocketConfig.fir@197383.4]
  assign _T_1459 = io_pmp_0_cfg_a[0] & _T_1457; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@197385.4]
  assign _T_1460 = io_pmp_0_cfg_a[1] ? _T_1401 : _T_1459; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@197386.4]
  assign _T_1461 = ~io_pmp_0_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@197387.4]
  assign _T_1462 = default_ & _T_1461; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@197388.4]
  assign _T_1500 = _T_1215[2:0] & _T_51; // @[PMP.scala 126:113:chipyard.TestHarness.RocketConfig.fir@197426.4]
  assign _T_1501 = _T_1500 != 3'h0; // @[PMP.scala 126:146:chipyard.TestHarness.RocketConfig.fir@197427.4]
  assign _T_1502 = _T_1225 & _T_1501; // @[PMP.scala 126:83:chipyard.TestHarness.RocketConfig.fir@197428.4]
  assign _T_1504 = ~_T_1502; // @[PMP.scala 127:24:chipyard.TestHarness.RocketConfig.fir@197430.4]
  assign _T_1506 = ~io_pmp_0_mask[2:0]; // @[PMP.scala 128:34:chipyard.TestHarness.RocketConfig.fir@197432.4]
  assign _T_1507 = _T_5 & _T_1506; // @[PMP.scala 128:32:chipyard.TestHarness.RocketConfig.fir@197433.4]
  assign _T_1508 = _T_1507 == 3'h0; // @[PMP.scala 128:57:chipyard.TestHarness.RocketConfig.fir@197434.4]
  assign _T_1510 = io_pmp_0_cfg_a[1] ? _T_1508 : _T_1504; // @[PMP.scala 129:8:chipyard.TestHarness.RocketConfig.fir@197436.4]
  assign _T_1562 = io_pmp_0_cfg_r | _T_1462; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@197496.4]
  assign _T_1563 = _T_1510 & _T_1562; // @[PMP.scala 183:26:chipyard.TestHarness.RocketConfig.fir@197497.4]
  assign _T_1564 = io_pmp_0_cfg_w | _T_1462; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@197499.4]
  assign _T_1565 = _T_1510 & _T_1564; // @[PMP.scala 184:26:chipyard.TestHarness.RocketConfig.fir@197500.4]
  assign _T_1566 = io_pmp_0_cfg_x | _T_1462; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@197502.4]
  assign _T_1567 = _T_1510 & _T_1566; // @[PMP.scala 185:26:chipyard.TestHarness.RocketConfig.fir@197503.4]
  assign io_r = _T_1460 ? _T_1563 : _T_1372_cfg_r; // @[PMP.scala 189:8:chipyard.TestHarness.RocketConfig.fir@197506.4]
  assign io_w = _T_1460 ? _T_1565 : _T_1372_cfg_w; // @[PMP.scala 190:8:chipyard.TestHarness.RocketConfig.fir@197507.4]
  assign io_x = _T_1460 ? _T_1567 : _T_1372_cfg_x; // @[PMP.scala 191:8:chipyard.TestHarness.RocketConfig.fir@197508.4]
endmodule
