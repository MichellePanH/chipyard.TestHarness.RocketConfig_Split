module RoundAnyRawFNToRecFN_2( // @[:chipyard.TestHarness.RocketConfig.fir@235580.2]
  input         io_in_isZero, // @[:chipyard.TestHarness.RocketConfig.fir@235581.4]
  input         io_in_sign, // @[:chipyard.TestHarness.RocketConfig.fir@235581.4]
  input  [8:0]  io_in_sExp, // @[:chipyard.TestHarness.RocketConfig.fir@235581.4]
  input  [64:0] io_in_sig, // @[:chipyard.TestHarness.RocketConfig.fir@235581.4]
  input  [2:0]  io_roundingMode, // @[:chipyard.TestHarness.RocketConfig.fir@235581.4]
  output [64:0] io_out, // @[:chipyard.TestHarness.RocketConfig.fir@235581.4]
  output [4:0]  io_exceptionFlags // @[:chipyard.TestHarness.RocketConfig.fir@235581.4]
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53:chipyard.TestHarness.RocketConfig.fir@235584.4]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53:chipyard.TestHarness.RocketConfig.fir@235586.4]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53:chipyard.TestHarness.RocketConfig.fir@235587.4]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53:chipyard.TestHarness.RocketConfig.fir@235588.4]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53:chipyard.TestHarness.RocketConfig.fir@235589.4]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27:chipyard.TestHarness.RocketConfig.fir@235590.4]
  wire  _T_1; // @[RoundAnyRawFNToRecFN.scala 96:66:chipyard.TestHarness.RocketConfig.fir@235591.4]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63:chipyard.TestHarness.RocketConfig.fir@235592.4]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42:chipyard.TestHarness.RocketConfig.fir@235593.4]
  wire [11:0] _GEN_0; // @[RoundAnyRawFNToRecFN.scala 102:25:chipyard.TestHarness.RocketConfig.fir@235594.4]
  wire [12:0] _T_3; // @[RoundAnyRawFNToRecFN.scala 102:25:chipyard.TestHarness.RocketConfig.fir@235594.4]
  wire [12:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 104:31:chipyard.TestHarness.RocketConfig.fir@235596.4]
  wire  _T_7; // @[RoundAnyRawFNToRecFN.scala 115:60:chipyard.TestHarness.RocketConfig.fir@235599.4]
  wire [55:0] adjustedSig; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@235600.4]
  wire [55:0] _T_14; // @[RoundAnyRawFNToRecFN.scala 162:40:chipyard.TestHarness.RocketConfig.fir@235619.4]
  wire  _T_15; // @[RoundAnyRawFNToRecFN.scala 162:56:chipyard.TestHarness.RocketConfig.fir@235620.4]
  wire [55:0] _T_16; // @[RoundAnyRawFNToRecFN.scala 163:42:chipyard.TestHarness.RocketConfig.fir@235621.4]
  wire  _T_17; // @[RoundAnyRawFNToRecFN.scala 163:62:chipyard.TestHarness.RocketConfig.fir@235622.4]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 164:36:chipyard.TestHarness.RocketConfig.fir@235623.4]
  wire  _T_19; // @[RoundAnyRawFNToRecFN.scala 167:38:chipyard.TestHarness.RocketConfig.fir@235624.4]
  wire  _T_20; // @[RoundAnyRawFNToRecFN.scala 167:67:chipyard.TestHarness.RocketConfig.fir@235625.4]
  wire  _T_21; // @[RoundAnyRawFNToRecFN.scala 169:29:chipyard.TestHarness.RocketConfig.fir@235626.4]
  wire  _T_22; // @[RoundAnyRawFNToRecFN.scala 168:31:chipyard.TestHarness.RocketConfig.fir@235627.4]
  wire [55:0] _T_23; // @[RoundAnyRawFNToRecFN.scala 172:32:chipyard.TestHarness.RocketConfig.fir@235628.4]
  wire [54:0] _T_25; // @[RoundAnyRawFNToRecFN.scala 172:49:chipyard.TestHarness.RocketConfig.fir@235630.4]
  wire  _T_26; // @[RoundAnyRawFNToRecFN.scala 173:49:chipyard.TestHarness.RocketConfig.fir@235631.4]
  wire  _T_27; // @[RoundAnyRawFNToRecFN.scala 174:30:chipyard.TestHarness.RocketConfig.fir@235632.4]
  wire  _T_28; // @[RoundAnyRawFNToRecFN.scala 173:64:chipyard.TestHarness.RocketConfig.fir@235633.4]
  wire [54:0] _T_30; // @[RoundAnyRawFNToRecFN.scala 173:25:chipyard.TestHarness.RocketConfig.fir@235635.4]
  wire [54:0] _T_31; // @[RoundAnyRawFNToRecFN.scala 173:21:chipyard.TestHarness.RocketConfig.fir@235636.4]
  wire [54:0] _T_32; // @[RoundAnyRawFNToRecFN.scala 172:61:chipyard.TestHarness.RocketConfig.fir@235637.4]
  wire [55:0] _T_34; // @[RoundAnyRawFNToRecFN.scala 178:30:chipyard.TestHarness.RocketConfig.fir@235639.4]
  wire  _T_36; // @[RoundAnyRawFNToRecFN.scala 179:42:chipyard.TestHarness.RocketConfig.fir@235641.4]
  wire [54:0] _T_38; // @[RoundAnyRawFNToRecFN.scala 179:24:chipyard.TestHarness.RocketConfig.fir@235643.4]
  wire [54:0] _GEN_1; // @[RoundAnyRawFNToRecFN.scala 178:47:chipyard.TestHarness.RocketConfig.fir@235644.4]
  wire [54:0] _T_39; // @[RoundAnyRawFNToRecFN.scala 178:47:chipyard.TestHarness.RocketConfig.fir@235644.4]
  wire [54:0] _T_40; // @[RoundAnyRawFNToRecFN.scala 171:16:chipyard.TestHarness.RocketConfig.fir@235645.4]
  wire [2:0] _T_42; // @[RoundAnyRawFNToRecFN.scala 183:69:chipyard.TestHarness.RocketConfig.fir@235647.4]
  wire [12:0] _GEN_2; // @[RoundAnyRawFNToRecFN.scala 183:40:chipyard.TestHarness.RocketConfig.fir@235648.4]
  wire [13:0] _T_43; // @[RoundAnyRawFNToRecFN.scala 183:40:chipyard.TestHarness.RocketConfig.fir@235648.4]
  wire [11:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37:chipyard.TestHarness.RocketConfig.fir@235649.4]
  wire [51:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 189:27:chipyard.TestHarness.RocketConfig.fir@235652.4]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:64:chipyard.TestHarness.RocketConfig.fir@235680.4]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:43:chipyard.TestHarness.RocketConfig.fir@235684.4]
  wire [11:0] _T_75; // @[RoundAnyRawFNToRecFN.scala 251:18:chipyard.TestHarness.RocketConfig.fir@235697.4]
  wire [11:0] _T_76; // @[RoundAnyRawFNToRecFN.scala 251:14:chipyard.TestHarness.RocketConfig.fir@235698.4]
  wire [11:0] expOut; // @[RoundAnyRawFNToRecFN.scala 250:24:chipyard.TestHarness.RocketConfig.fir@235699.4]
  wire [51:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12:chipyard.TestHarness.RocketConfig.fir@235721.4]
  wire [12:0] _T_101; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@235725.4]
  wire [1:0] _T_103; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@235728.4]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53:chipyard.TestHarness.RocketConfig.fir@235584.4]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53:chipyard.TestHarness.RocketConfig.fir@235586.4]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53:chipyard.TestHarness.RocketConfig.fir@235587.4]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53:chipyard.TestHarness.RocketConfig.fir@235588.4]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53:chipyard.TestHarness.RocketConfig.fir@235589.4]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27:chipyard.TestHarness.RocketConfig.fir@235590.4]
  assign _T_1 = ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:66:chipyard.TestHarness.RocketConfig.fir@235591.4]
  assign _T_2 = roundingMode_max & _T_1; // @[RoundAnyRawFNToRecFN.scala 96:63:chipyard.TestHarness.RocketConfig.fir@235592.4]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42:chipyard.TestHarness.RocketConfig.fir@235593.4]
  assign _GEN_0 = {{3{io_in_sExp[8]}},io_in_sExp}; // @[RoundAnyRawFNToRecFN.scala 102:25:chipyard.TestHarness.RocketConfig.fir@235594.4]
  assign _T_3 = $signed(_GEN_0) + 12'sh780; // @[RoundAnyRawFNToRecFN.scala 102:25:chipyard.TestHarness.RocketConfig.fir@235594.4]
  assign sAdjustedExp = {1'b0,$signed(_T_3[11:0])}; // @[RoundAnyRawFNToRecFN.scala 104:31:chipyard.TestHarness.RocketConfig.fir@235596.4]
  assign _T_7 = |io_in_sig[9:0]; // @[RoundAnyRawFNToRecFN.scala 115:60:chipyard.TestHarness.RocketConfig.fir@235599.4]
  assign adjustedSig = {io_in_sig[64:10],_T_7}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@235600.4]
  assign _T_14 = adjustedSig & 56'h2; // @[RoundAnyRawFNToRecFN.scala 162:40:chipyard.TestHarness.RocketConfig.fir@235619.4]
  assign _T_15 = |_T_14; // @[RoundAnyRawFNToRecFN.scala 162:56:chipyard.TestHarness.RocketConfig.fir@235620.4]
  assign _T_16 = adjustedSig & 56'h1; // @[RoundAnyRawFNToRecFN.scala 163:42:chipyard.TestHarness.RocketConfig.fir@235621.4]
  assign _T_17 = |_T_16; // @[RoundAnyRawFNToRecFN.scala 163:62:chipyard.TestHarness.RocketConfig.fir@235622.4]
  assign common_inexact = _T_15 | _T_17; // @[RoundAnyRawFNToRecFN.scala 164:36:chipyard.TestHarness.RocketConfig.fir@235623.4]
  assign _T_19 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38:chipyard.TestHarness.RocketConfig.fir@235624.4]
  assign _T_20 = _T_19 & _T_15; // @[RoundAnyRawFNToRecFN.scala 167:67:chipyard.TestHarness.RocketConfig.fir@235625.4]
  assign _T_21 = roundMagUp & common_inexact; // @[RoundAnyRawFNToRecFN.scala 169:29:chipyard.TestHarness.RocketConfig.fir@235626.4]
  assign _T_22 = _T_20 | _T_21; // @[RoundAnyRawFNToRecFN.scala 168:31:chipyard.TestHarness.RocketConfig.fir@235627.4]
  assign _T_23 = adjustedSig | 56'h3; // @[RoundAnyRawFNToRecFN.scala 172:32:chipyard.TestHarness.RocketConfig.fir@235628.4]
  assign _T_25 = _T_23[55:2] + 54'h1; // @[RoundAnyRawFNToRecFN.scala 172:49:chipyard.TestHarness.RocketConfig.fir@235630.4]
  assign _T_26 = roundingMode_near_even & _T_15; // @[RoundAnyRawFNToRecFN.scala 173:49:chipyard.TestHarness.RocketConfig.fir@235631.4]
  assign _T_27 = ~_T_17; // @[RoundAnyRawFNToRecFN.scala 174:30:chipyard.TestHarness.RocketConfig.fir@235632.4]
  assign _T_28 = _T_26 & _T_27; // @[RoundAnyRawFNToRecFN.scala 173:64:chipyard.TestHarness.RocketConfig.fir@235633.4]
  assign _T_30 = _T_28 ? 55'h1 : 55'h0; // @[RoundAnyRawFNToRecFN.scala 173:25:chipyard.TestHarness.RocketConfig.fir@235635.4]
  assign _T_31 = ~_T_30; // @[RoundAnyRawFNToRecFN.scala 173:21:chipyard.TestHarness.RocketConfig.fir@235636.4]
  assign _T_32 = _T_25 & _T_31; // @[RoundAnyRawFNToRecFN.scala 172:61:chipyard.TestHarness.RocketConfig.fir@235637.4]
  assign _T_34 = adjustedSig & 56'hfffffffffffffc; // @[RoundAnyRawFNToRecFN.scala 178:30:chipyard.TestHarness.RocketConfig.fir@235639.4]
  assign _T_36 = roundingMode_odd & common_inexact; // @[RoundAnyRawFNToRecFN.scala 179:42:chipyard.TestHarness.RocketConfig.fir@235641.4]
  assign _T_38 = _T_36 ? 55'h1 : 55'h0; // @[RoundAnyRawFNToRecFN.scala 179:24:chipyard.TestHarness.RocketConfig.fir@235643.4]
  assign _GEN_1 = {{1'd0}, _T_34[55:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47:chipyard.TestHarness.RocketConfig.fir@235644.4]
  assign _T_39 = _GEN_1 | _T_38; // @[RoundAnyRawFNToRecFN.scala 178:47:chipyard.TestHarness.RocketConfig.fir@235644.4]
  assign _T_40 = _T_22 ? _T_32 : _T_39; // @[RoundAnyRawFNToRecFN.scala 171:16:chipyard.TestHarness.RocketConfig.fir@235645.4]
  assign _T_42 = {1'b0,$signed(_T_40[54:53])}; // @[RoundAnyRawFNToRecFN.scala 183:69:chipyard.TestHarness.RocketConfig.fir@235647.4]
  assign _GEN_2 = {{10{_T_42[2]}},_T_42}; // @[RoundAnyRawFNToRecFN.scala 183:40:chipyard.TestHarness.RocketConfig.fir@235648.4]
  assign _T_43 = $signed(sAdjustedExp) + $signed(_GEN_2); // @[RoundAnyRawFNToRecFN.scala 183:40:chipyard.TestHarness.RocketConfig.fir@235648.4]
  assign common_expOut = _T_43[11:0]; // @[RoundAnyRawFNToRecFN.scala 185:37:chipyard.TestHarness.RocketConfig.fir@235649.4]
  assign common_fractOut = _T_40[51:0]; // @[RoundAnyRawFNToRecFN.scala 189:27:chipyard.TestHarness.RocketConfig.fir@235652.4]
  assign commonCase = ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:64:chipyard.TestHarness.RocketConfig.fir@235680.4]
  assign inexact = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43:chipyard.TestHarness.RocketConfig.fir@235684.4]
  assign _T_75 = io_in_isZero ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18:chipyard.TestHarness.RocketConfig.fir@235697.4]
  assign _T_76 = ~_T_75; // @[RoundAnyRawFNToRecFN.scala 251:14:chipyard.TestHarness.RocketConfig.fir@235698.4]
  assign expOut = common_expOut & _T_76; // @[RoundAnyRawFNToRecFN.scala 250:24:chipyard.TestHarness.RocketConfig.fir@235699.4]
  assign fractOut = io_in_isZero ? 52'h0 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12:chipyard.TestHarness.RocketConfig.fir@235721.4]
  assign _T_101 = {io_in_sign,expOut}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@235725.4]
  assign _T_103 = {1'h0,inexact}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@235728.4]
  assign io_out = {_T_101,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12:chipyard.TestHarness.RocketConfig.fir@235727.4]
  assign io_exceptionFlags = {3'h0,_T_103}; // @[RoundAnyRawFNToRecFN.scala 285:23:chipyard.TestHarness.RocketConfig.fir@235732.4]
endmodule
