module DCacheModuleImpl_Anon_2( // @[:chipyard.TestHarness.RocketConfig.fir@213738.2]
  input         io_in_0_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [11:0] io_in_0_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input         io_in_0_bits_write, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [63:0] io_in_0_bits_wdata, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [7:0]  io_in_0_bits_eccMask, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [3:0]  io_in_0_bits_way_en, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  output        io_in_1_ready, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input         io_in_1_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [11:0] io_in_1_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input         io_in_1_bits_write, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [63:0] io_in_1_bits_wdata, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [7:0]  io_in_1_bits_eccMask, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [3:0]  io_in_1_bits_way_en, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  output        io_in_2_ready, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input         io_in_2_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [11:0] io_in_2_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [63:0] io_in_2_bits_wdata, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [7:0]  io_in_2_bits_eccMask, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  output        io_in_3_ready, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input         io_in_3_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [11:0] io_in_3_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [63:0] io_in_3_bits_wdata, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  input  [7:0]  io_in_3_bits_eccMask, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  output        io_out_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  output [11:0] io_out_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  output        io_out_bits_write, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  output [63:0] io_out_bits_wdata, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  output [7:0]  io_out_bits_eccMask, // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
  output [3:0]  io_out_bits_way_en // @[:chipyard.TestHarness.RocketConfig.fir@213741.4]
);
  wire [7:0] _GEN_2; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213750.4]
  wire [63:0] _GEN_4; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213750.4]
  wire [11:0] _GEN_6; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213750.4]
  wire [3:0] _GEN_8; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213759.4]
  wire [7:0] _GEN_9; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213759.4]
  wire [63:0] _GEN_11; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213759.4]
  wire  _GEN_12; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213759.4]
  wire [11:0] _GEN_13; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213759.4]
  wire  _T; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213777.4]
  wire  _T_1; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213778.4]
  wire  grant_3; // @[Arbiter.scala 31:78:chipyard.TestHarness.RocketConfig.fir@213781.4]
  wire  _T_6; // @[Arbiter.scala 135:19:chipyard.TestHarness.RocketConfig.fir@213790.4]
  assign _GEN_2 = io_in_2_valid ? io_in_2_bits_eccMask : io_in_3_bits_eccMask; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213750.4]
  assign _GEN_4 = io_in_2_valid ? io_in_2_bits_wdata : io_in_3_bits_wdata; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213750.4]
  assign _GEN_6 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213750.4]
  assign _GEN_8 = io_in_1_valid ? io_in_1_bits_way_en : 4'hf; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213759.4]
  assign _GEN_9 = io_in_1_valid ? 8'hff : _GEN_2; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213759.4]
  assign _GEN_11 = io_in_1_valid ? io_in_1_bits_wdata : _GEN_4; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213759.4]
  assign _GEN_12 = io_in_1_valid & io_in_1_bits_write; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213759.4]
  assign _GEN_13 = io_in_1_valid ? io_in_1_bits_addr : _GEN_6; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213759.4]
  assign _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213777.4]
  assign _T_1 = _T | io_in_2_valid; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213778.4]
  assign grant_3 = ~_T_1; // @[Arbiter.scala 31:78:chipyard.TestHarness.RocketConfig.fir@213781.4]
  assign _T_6 = ~grant_3; // @[Arbiter.scala 135:19:chipyard.TestHarness.RocketConfig.fir@213790.4]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 134:14:chipyard.TestHarness.RocketConfig.fir@213785.4]
  assign io_in_2_ready = ~_T; // @[Arbiter.scala 134:14:chipyard.TestHarness.RocketConfig.fir@213787.4]
  assign io_in_3_ready = ~_T_1; // @[Arbiter.scala 134:14:chipyard.TestHarness.RocketConfig.fir@213789.4]
  assign io_out_valid = _T_6 | io_in_3_valid; // @[Arbiter.scala 135:16:chipyard.TestHarness.RocketConfig.fir@213792.4]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_13; // @[Arbiter.scala 124:15:chipyard.TestHarness.RocketConfig.fir@213749.4 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213757.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213766.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213775.6]
  assign io_out_bits_write = io_in_0_valid ? io_in_0_bits_write : _GEN_12; // @[Arbiter.scala 124:15:chipyard.TestHarness.RocketConfig.fir@213748.4 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213756.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213765.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213774.6]
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : _GEN_11; // @[Arbiter.scala 124:15:chipyard.TestHarness.RocketConfig.fir@213747.4 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213755.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213764.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213773.6]
  assign io_out_bits_eccMask = io_in_0_valid ? io_in_0_bits_eccMask : _GEN_9; // @[Arbiter.scala 124:15:chipyard.TestHarness.RocketConfig.fir@213745.4 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213753.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213762.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213771.6]
  assign io_out_bits_way_en = io_in_0_valid ? io_in_0_bits_way_en : _GEN_8; // @[Arbiter.scala 124:15:chipyard.TestHarness.RocketConfig.fir@213744.4 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213752.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213761.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213770.6]
endmodule
