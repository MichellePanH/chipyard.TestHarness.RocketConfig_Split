module IntSyncSyncCrossingSink_1( // @[:chipyard.TestHarness.RocketConfig.fir@233304.2]
  input   auto_in_sync_0, // @[:chipyard.TestHarness.RocketConfig.fir@233307.4]
  output  auto_out_0 // @[:chipyard.TestHarness.RocketConfig.fir@233307.4]
);
  assign auto_out_0 = auto_in_sync_0; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@233316.4]
endmodule
