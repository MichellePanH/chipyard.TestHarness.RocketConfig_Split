module Atomics( // @[:chipyard.TestHarness.RocketConfig.fir@84623.2]
  input         io_write, // @[:chipyard.TestHarness.RocketConfig.fir@84626.4]
  input  [2:0]  io_a_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@84626.4]
  input  [2:0]  io_a_param, // @[:chipyard.TestHarness.RocketConfig.fir@84626.4]
  input  [7:0]  io_a_mask, // @[:chipyard.TestHarness.RocketConfig.fir@84626.4]
  input  [63:0] io_a_data, // @[:chipyard.TestHarness.RocketConfig.fir@84626.4]
  input  [63:0] io_data_in, // @[:chipyard.TestHarness.RocketConfig.fir@84626.4]
  output [63:0] io_data_out // @[:chipyard.TestHarness.RocketConfig.fir@84626.4]
);
  wire  adder; // @[Atomics.scala 21:28:chipyard.TestHarness.RocketConfig.fir@84631.4]
  wire  unsigned_; // @[Atomics.scala 22:28:chipyard.TestHarness.RocketConfig.fir@84632.4]
  wire  take_max; // @[Atomics.scala 23:28:chipyard.TestHarness.RocketConfig.fir@84633.4]
  wire [7:0] _T; // @[Atomics.scala 25:42:chipyard.TestHarness.RocketConfig.fir@84634.4]
  wire [7:0] _T_2; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@84636.4]
  wire [7:0] signBit; // @[Atomics.scala 25:27:chipyard.TestHarness.RocketConfig.fir@84637.4]
  wire [63:0] _T_3; // @[Atomics.scala 26:38:chipyard.TestHarness.RocketConfig.fir@84638.4]
  wire [63:0] inv_d; // @[Atomics.scala 26:18:chipyard.TestHarness.RocketConfig.fir@84639.4]
  wire [7:0] _T_13; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84649.4]
  wire [7:0] _T_15; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84651.4]
  wire [7:0] _T_17; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84653.4]
  wire [7:0] _T_19; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84655.4]
  wire [7:0] _T_21; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84657.4]
  wire [7:0] _T_23; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84659.4]
  wire [7:0] _T_25; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84661.4]
  wire [7:0] _T_27; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84663.4]
  wire [63:0] _T_34; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@84670.4]
  wire [63:0] _T_35; // @[Atomics.scala 27:44:chipyard.TestHarness.RocketConfig.fir@84671.4]
  wire [63:0] sum; // @[Atomics.scala 27:57:chipyard.TestHarness.RocketConfig.fir@84673.4]
  wire [7:0] _T_107; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@84744.4]
  wire [7:0] _T_108; // @[Atomics.scala 28:83:chipyard.TestHarness.RocketConfig.fir@84745.4]
  wire  sign_a; // @[Atomics.scala 28:97:chipyard.TestHarness.RocketConfig.fir@84746.4]
  wire [7:0] _T_179; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@84817.4]
  wire [7:0] _T_180; // @[Atomics.scala 28:83:chipyard.TestHarness.RocketConfig.fir@84818.4]
  wire  sign_d; // @[Atomics.scala 28:97:chipyard.TestHarness.RocketConfig.fir@84819.4]
  wire [7:0] _T_251; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@84890.4]
  wire [7:0] _T_252; // @[Atomics.scala 28:83:chipyard.TestHarness.RocketConfig.fir@84891.4]
  wire  sign_s; // @[Atomics.scala 28:97:chipyard.TestHarness.RocketConfig.fir@84892.4]
  wire  a_bigger_uneq; // @[Atomics.scala 32:32:chipyard.TestHarness.RocketConfig.fir@84893.4]
  wire  _T_253; // @[Atomics.scala 33:29:chipyard.TestHarness.RocketConfig.fir@84894.4]
  wire  _T_254; // @[Atomics.scala 33:41:chipyard.TestHarness.RocketConfig.fir@84895.4]
  wire  a_bigger; // @[Atomics.scala 33:21:chipyard.TestHarness.RocketConfig.fir@84896.4]
  wire  pick_a; // @[Atomics.scala 34:25:chipyard.TestHarness.RocketConfig.fir@84897.4]
  wire [1:0] _T_385; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85033.4]
  wire [3:0] _GEN_1; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85034.4]
  wire [3:0] _GEN_2; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85034.4]
  wire [3:0] _GEN_3; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85034.4]
  wire [3:0] _T_386; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85034.4]
  wire [1:0] _T_388; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85036.4]
  wire [3:0] _T_389; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85037.4]
  wire [1:0] _T_391; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85039.4]
  wire [3:0] _T_392; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85040.4]
  wire [1:0] _T_394; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85042.4]
  wire [3:0] _T_395; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85043.4]
  wire [1:0] _T_397; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85045.4]
  wire [3:0] _T_398; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85046.4]
  wire [1:0] _T_400; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85048.4]
  wire [3:0] _T_401; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85049.4]
  wire [1:0] _T_403; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85051.4]
  wire [3:0] _T_404; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85052.4]
  wire [1:0] _T_406; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85054.4]
  wire [3:0] _T_407; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85055.4]
  wire [1:0] _T_409; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85057.4]
  wire [3:0] _T_410; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85058.4]
  wire [1:0] _T_412; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85060.4]
  wire [3:0] _T_413; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85061.4]
  wire [1:0] _T_415; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85063.4]
  wire [3:0] _T_416; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85064.4]
  wire [1:0] _T_418; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85066.4]
  wire [3:0] _T_419; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85067.4]
  wire [1:0] _T_421; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85069.4]
  wire [3:0] _T_422; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85070.4]
  wire [1:0] _T_424; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85072.4]
  wire [3:0] _T_425; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85073.4]
  wire [1:0] _T_427; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85075.4]
  wire [3:0] _T_428; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85076.4]
  wire [1:0] _T_430; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85078.4]
  wire [3:0] _T_431; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85079.4]
  wire [1:0] _T_433; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85081.4]
  wire [3:0] _T_434; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85082.4]
  wire [1:0] _T_436; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85084.4]
  wire [3:0] _T_437; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85085.4]
  wire [1:0] _T_439; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85087.4]
  wire [3:0] _T_440; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85088.4]
  wire [1:0] _T_442; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85090.4]
  wire [3:0] _T_443; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85091.4]
  wire [1:0] _T_445; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85093.4]
  wire [3:0] _T_446; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85094.4]
  wire [1:0] _T_448; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85096.4]
  wire [3:0] _T_449; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85097.4]
  wire [1:0] _T_451; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85099.4]
  wire [3:0] _T_452; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85100.4]
  wire [1:0] _T_454; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85102.4]
  wire [3:0] _T_455; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85103.4]
  wire [1:0] _T_457; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85105.4]
  wire [3:0] _T_458; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85106.4]
  wire [1:0] _T_460; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85108.4]
  wire [3:0] _T_461; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85109.4]
  wire [1:0] _T_463; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85111.4]
  wire [3:0] _T_464; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85112.4]
  wire [1:0] _T_466; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85114.4]
  wire [3:0] _T_467; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85115.4]
  wire [1:0] _T_469; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85117.4]
  wire [3:0] _T_470; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85118.4]
  wire [1:0] _T_472; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85120.4]
  wire [3:0] _T_473; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85121.4]
  wire [1:0] _T_475; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85123.4]
  wire [3:0] _T_476; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85124.4]
  wire [1:0] _T_478; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85126.4]
  wire [3:0] _T_479; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85127.4]
  wire [1:0] _T_481; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85129.4]
  wire [3:0] _T_482; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85130.4]
  wire [1:0] _T_484; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85132.4]
  wire [3:0] _T_485; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85133.4]
  wire [1:0] _T_487; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85135.4]
  wire [3:0] _T_488; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85136.4]
  wire [1:0] _T_490; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85138.4]
  wire [3:0] _T_491; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85139.4]
  wire [1:0] _T_493; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85141.4]
  wire [3:0] _T_494; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85142.4]
  wire [1:0] _T_496; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85144.4]
  wire [3:0] _T_497; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85145.4]
  wire [1:0] _T_499; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85147.4]
  wire [3:0] _T_500; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85148.4]
  wire [1:0] _T_502; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85150.4]
  wire [3:0] _T_503; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85151.4]
  wire [1:0] _T_505; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85153.4]
  wire [3:0] _T_506; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85154.4]
  wire [1:0] _T_508; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85156.4]
  wire [3:0] _T_509; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85157.4]
  wire [1:0] _T_511; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85159.4]
  wire [3:0] _T_512; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85160.4]
  wire [1:0] _T_514; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85162.4]
  wire [3:0] _T_515; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85163.4]
  wire [1:0] _T_517; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85165.4]
  wire [3:0] _T_518; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85166.4]
  wire [1:0] _T_520; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85168.4]
  wire [3:0] _T_521; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85169.4]
  wire [1:0] _T_523; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85171.4]
  wire [3:0] _T_524; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85172.4]
  wire [1:0] _T_526; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85174.4]
  wire [3:0] _T_527; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85175.4]
  wire [1:0] _T_529; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85177.4]
  wire [3:0] _T_530; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85178.4]
  wire [1:0] _T_532; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85180.4]
  wire [3:0] _T_533; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85181.4]
  wire [1:0] _T_535; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85183.4]
  wire [3:0] _T_536; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85184.4]
  wire [1:0] _T_538; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85186.4]
  wire [3:0] _T_539; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85187.4]
  wire [1:0] _T_541; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85189.4]
  wire [3:0] _T_542; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85190.4]
  wire [1:0] _T_544; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85192.4]
  wire [3:0] _T_545; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85193.4]
  wire [1:0] _T_547; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85195.4]
  wire [3:0] _T_548; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85196.4]
  wire [1:0] _T_550; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85198.4]
  wire [3:0] _T_551; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85199.4]
  wire [1:0] _T_553; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85201.4]
  wire [3:0] _T_554; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85202.4]
  wire [1:0] _T_556; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85204.4]
  wire [3:0] _T_557; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85205.4]
  wire [1:0] _T_559; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85207.4]
  wire [3:0] _T_560; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85208.4]
  wire [1:0] _T_562; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85210.4]
  wire [3:0] _T_563; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85211.4]
  wire [1:0] _T_565; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85213.4]
  wire [3:0] _T_566; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85214.4]
  wire [1:0] _T_568; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85216.4]
  wire [3:0] _T_569; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85217.4]
  wire [1:0] _T_571; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85219.4]
  wire [3:0] _T_572; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85220.4]
  wire [1:0] _T_574; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85222.4]
  wire [3:0] _T_575; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85223.4]
  wire [7:0] _T_583; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85231.4]
  wire [15:0] _T_591; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85239.4]
  wire [7:0] _T_598; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85246.4]
  wire [31:0] _T_607; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85255.4]
  wire [7:0] _T_614; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85262.4]
  wire [15:0] _T_622; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85270.4]
  wire [7:0] _T_629; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85277.4]
  wire [31:0] _T_638; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85286.4]
  wire [63:0] logical; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85287.4]
  wire [1:0] _T_640; // @[Atomics.scala 51:8:chipyard.TestHarness.RocketConfig.fir@85289.4]
  wire [1:0] _GEN_6; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  wire [1:0] _GEN_7; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  wire [1:0] _GEN_8; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  wire [1:0] _GEN_9; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  wire [1:0] _GEN_10; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  wire [1:0] _GEN_11; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  wire [1:0] select; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  wire [1:0] selects_0; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85309.4]
  wire [1:0] selects_1; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85310.4]
  wire [1:0] selects_2; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85311.4]
  wire [1:0] selects_3; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85312.4]
  wire [1:0] selects_4; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85313.4]
  wire [1:0] selects_5; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85314.4]
  wire [1:0] selects_6; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85315.4]
  wire [1:0] selects_7; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85316.4]
  wire [7:0] _GEN_13; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85397.4]
  wire [7:0] _GEN_14; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85397.4]
  wire [7:0] _GEN_15; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85397.4]
  wire [7:0] _GEN_17; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85397.4]
  wire [7:0] _GEN_18; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85397.4]
  wire [7:0] _GEN_19; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85397.4]
  wire [7:0] _GEN_21; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85398.4]
  wire [7:0] _GEN_22; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85398.4]
  wire [7:0] _GEN_23; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85398.4]
  wire [7:0] _GEN_25; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85398.4]
  wire [7:0] _GEN_26; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85398.4]
  wire [7:0] _GEN_27; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85398.4]
  wire [31:0] _T_692; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85399.4]
  wire [7:0] _GEN_29; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85400.4]
  wire [7:0] _GEN_30; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85400.4]
  wire [7:0] _GEN_31; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85400.4]
  wire [7:0] _GEN_33; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85400.4]
  wire [7:0] _GEN_34; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85400.4]
  wire [7:0] _GEN_35; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85400.4]
  wire [7:0] _GEN_37; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85401.4]
  wire [7:0] _GEN_38; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85401.4]
  wire [7:0] _GEN_39; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85401.4]
  wire [7:0] _GEN_41; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85401.4]
  wire [7:0] _GEN_42; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85401.4]
  wire [7:0] _GEN_43; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85401.4]
  wire [31:0] _T_695; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85402.4]
  assign adder = io_a_param[2]; // @[Atomics.scala 21:28:chipyard.TestHarness.RocketConfig.fir@84631.4]
  assign unsigned_ = io_a_param[1]; // @[Atomics.scala 22:28:chipyard.TestHarness.RocketConfig.fir@84632.4]
  assign take_max = io_a_param[0]; // @[Atomics.scala 23:28:chipyard.TestHarness.RocketConfig.fir@84633.4]
  assign _T = ~io_a_mask; // @[Atomics.scala 25:42:chipyard.TestHarness.RocketConfig.fir@84634.4]
  assign _T_2 = {1'h1,_T[7:1]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@84636.4]
  assign signBit = io_a_mask & _T_2; // @[Atomics.scala 25:27:chipyard.TestHarness.RocketConfig.fir@84637.4]
  assign _T_3 = ~io_data_in; // @[Atomics.scala 26:38:chipyard.TestHarness.RocketConfig.fir@84638.4]
  assign inv_d = adder ? io_data_in : _T_3; // @[Atomics.scala 26:18:chipyard.TestHarness.RocketConfig.fir@84639.4]
  assign _T_13 = io_a_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84649.4]
  assign _T_15 = io_a_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84651.4]
  assign _T_17 = io_a_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84653.4]
  assign _T_19 = io_a_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84655.4]
  assign _T_21 = io_a_mask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84657.4]
  assign _T_23 = io_a_mask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84659.4]
  assign _T_25 = io_a_mask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84661.4]
  assign _T_27 = io_a_mask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@84663.4]
  assign _T_34 = {_T_27,_T_25,_T_23,_T_21,_T_19,_T_17,_T_15,_T_13}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@84670.4]
  assign _T_35 = _T_34 & io_a_data; // @[Atomics.scala 27:44:chipyard.TestHarness.RocketConfig.fir@84671.4]
  assign sum = _T_35 + inv_d; // @[Atomics.scala 27:57:chipyard.TestHarness.RocketConfig.fir@84673.4]
  assign _T_107 = {io_a_data[63],io_a_data[55],io_a_data[47],io_a_data[39],io_a_data[31],io_a_data[23],io_a_data[15],io_a_data[7]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@84744.4]
  assign _T_108 = _T_107 & signBit; // @[Atomics.scala 28:83:chipyard.TestHarness.RocketConfig.fir@84745.4]
  assign sign_a = |_T_108; // @[Atomics.scala 28:97:chipyard.TestHarness.RocketConfig.fir@84746.4]
  assign _T_179 = {io_data_in[63],io_data_in[55],io_data_in[47],io_data_in[39],io_data_in[31],io_data_in[23],io_data_in[15],io_data_in[7]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@84817.4]
  assign _T_180 = _T_179 & signBit; // @[Atomics.scala 28:83:chipyard.TestHarness.RocketConfig.fir@84818.4]
  assign sign_d = |_T_180; // @[Atomics.scala 28:97:chipyard.TestHarness.RocketConfig.fir@84819.4]
  assign _T_251 = {sum[63],sum[55],sum[47],sum[39],sum[31],sum[23],sum[15],sum[7]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@84890.4]
  assign _T_252 = _T_251 & signBit; // @[Atomics.scala 28:83:chipyard.TestHarness.RocketConfig.fir@84891.4]
  assign sign_s = |_T_252; // @[Atomics.scala 28:97:chipyard.TestHarness.RocketConfig.fir@84892.4]
  assign a_bigger_uneq = unsigned_ == sign_a; // @[Atomics.scala 32:32:chipyard.TestHarness.RocketConfig.fir@84893.4]
  assign _T_253 = sign_a == sign_d; // @[Atomics.scala 33:29:chipyard.TestHarness.RocketConfig.fir@84894.4]
  assign _T_254 = ~sign_s; // @[Atomics.scala 33:41:chipyard.TestHarness.RocketConfig.fir@84895.4]
  assign a_bigger = _T_253 ? _T_254 : a_bigger_uneq; // @[Atomics.scala 33:21:chipyard.TestHarness.RocketConfig.fir@84896.4]
  assign pick_a = take_max == a_bigger; // @[Atomics.scala 34:25:chipyard.TestHarness.RocketConfig.fir@84897.4]
  assign _T_385 = {io_a_data[0],io_data_in[0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85033.4]
  assign _GEN_1 = 2'h1 == io_a_param[1:0] ? 4'he : 4'h6; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85034.4]
  assign _GEN_2 = 2'h2 == io_a_param[1:0] ? 4'h8 : _GEN_1; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85034.4]
  assign _GEN_3 = 2'h3 == io_a_param[1:0] ? 4'hc : _GEN_2; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85034.4]
  assign _T_386 = _GEN_3 >> _T_385; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85034.4]
  assign _T_388 = {io_a_data[1],io_data_in[1]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85036.4]
  assign _T_389 = _GEN_3 >> _T_388; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85037.4]
  assign _T_391 = {io_a_data[2],io_data_in[2]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85039.4]
  assign _T_392 = _GEN_3 >> _T_391; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85040.4]
  assign _T_394 = {io_a_data[3],io_data_in[3]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85042.4]
  assign _T_395 = _GEN_3 >> _T_394; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85043.4]
  assign _T_397 = {io_a_data[4],io_data_in[4]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85045.4]
  assign _T_398 = _GEN_3 >> _T_397; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85046.4]
  assign _T_400 = {io_a_data[5],io_data_in[5]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85048.4]
  assign _T_401 = _GEN_3 >> _T_400; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85049.4]
  assign _T_403 = {io_a_data[6],io_data_in[6]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85051.4]
  assign _T_404 = _GEN_3 >> _T_403; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85052.4]
  assign _T_406 = {io_a_data[7],io_data_in[7]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85054.4]
  assign _T_407 = _GEN_3 >> _T_406; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85055.4]
  assign _T_409 = {io_a_data[8],io_data_in[8]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85057.4]
  assign _T_410 = _GEN_3 >> _T_409; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85058.4]
  assign _T_412 = {io_a_data[9],io_data_in[9]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85060.4]
  assign _T_413 = _GEN_3 >> _T_412; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85061.4]
  assign _T_415 = {io_a_data[10],io_data_in[10]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85063.4]
  assign _T_416 = _GEN_3 >> _T_415; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85064.4]
  assign _T_418 = {io_a_data[11],io_data_in[11]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85066.4]
  assign _T_419 = _GEN_3 >> _T_418; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85067.4]
  assign _T_421 = {io_a_data[12],io_data_in[12]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85069.4]
  assign _T_422 = _GEN_3 >> _T_421; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85070.4]
  assign _T_424 = {io_a_data[13],io_data_in[13]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85072.4]
  assign _T_425 = _GEN_3 >> _T_424; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85073.4]
  assign _T_427 = {io_a_data[14],io_data_in[14]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85075.4]
  assign _T_428 = _GEN_3 >> _T_427; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85076.4]
  assign _T_430 = {io_a_data[15],io_data_in[15]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85078.4]
  assign _T_431 = _GEN_3 >> _T_430; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85079.4]
  assign _T_433 = {io_a_data[16],io_data_in[16]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85081.4]
  assign _T_434 = _GEN_3 >> _T_433; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85082.4]
  assign _T_436 = {io_a_data[17],io_data_in[17]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85084.4]
  assign _T_437 = _GEN_3 >> _T_436; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85085.4]
  assign _T_439 = {io_a_data[18],io_data_in[18]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85087.4]
  assign _T_440 = _GEN_3 >> _T_439; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85088.4]
  assign _T_442 = {io_a_data[19],io_data_in[19]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85090.4]
  assign _T_443 = _GEN_3 >> _T_442; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85091.4]
  assign _T_445 = {io_a_data[20],io_data_in[20]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85093.4]
  assign _T_446 = _GEN_3 >> _T_445; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85094.4]
  assign _T_448 = {io_a_data[21],io_data_in[21]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85096.4]
  assign _T_449 = _GEN_3 >> _T_448; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85097.4]
  assign _T_451 = {io_a_data[22],io_data_in[22]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85099.4]
  assign _T_452 = _GEN_3 >> _T_451; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85100.4]
  assign _T_454 = {io_a_data[23],io_data_in[23]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85102.4]
  assign _T_455 = _GEN_3 >> _T_454; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85103.4]
  assign _T_457 = {io_a_data[24],io_data_in[24]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85105.4]
  assign _T_458 = _GEN_3 >> _T_457; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85106.4]
  assign _T_460 = {io_a_data[25],io_data_in[25]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85108.4]
  assign _T_461 = _GEN_3 >> _T_460; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85109.4]
  assign _T_463 = {io_a_data[26],io_data_in[26]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85111.4]
  assign _T_464 = _GEN_3 >> _T_463; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85112.4]
  assign _T_466 = {io_a_data[27],io_data_in[27]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85114.4]
  assign _T_467 = _GEN_3 >> _T_466; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85115.4]
  assign _T_469 = {io_a_data[28],io_data_in[28]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85117.4]
  assign _T_470 = _GEN_3 >> _T_469; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85118.4]
  assign _T_472 = {io_a_data[29],io_data_in[29]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85120.4]
  assign _T_473 = _GEN_3 >> _T_472; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85121.4]
  assign _T_475 = {io_a_data[30],io_data_in[30]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85123.4]
  assign _T_476 = _GEN_3 >> _T_475; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85124.4]
  assign _T_478 = {io_a_data[31],io_data_in[31]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85126.4]
  assign _T_479 = _GEN_3 >> _T_478; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85127.4]
  assign _T_481 = {io_a_data[32],io_data_in[32]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85129.4]
  assign _T_482 = _GEN_3 >> _T_481; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85130.4]
  assign _T_484 = {io_a_data[33],io_data_in[33]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85132.4]
  assign _T_485 = _GEN_3 >> _T_484; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85133.4]
  assign _T_487 = {io_a_data[34],io_data_in[34]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85135.4]
  assign _T_488 = _GEN_3 >> _T_487; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85136.4]
  assign _T_490 = {io_a_data[35],io_data_in[35]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85138.4]
  assign _T_491 = _GEN_3 >> _T_490; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85139.4]
  assign _T_493 = {io_a_data[36],io_data_in[36]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85141.4]
  assign _T_494 = _GEN_3 >> _T_493; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85142.4]
  assign _T_496 = {io_a_data[37],io_data_in[37]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85144.4]
  assign _T_497 = _GEN_3 >> _T_496; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85145.4]
  assign _T_499 = {io_a_data[38],io_data_in[38]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85147.4]
  assign _T_500 = _GEN_3 >> _T_499; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85148.4]
  assign _T_502 = {io_a_data[39],io_data_in[39]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85150.4]
  assign _T_503 = _GEN_3 >> _T_502; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85151.4]
  assign _T_505 = {io_a_data[40],io_data_in[40]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85153.4]
  assign _T_506 = _GEN_3 >> _T_505; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85154.4]
  assign _T_508 = {io_a_data[41],io_data_in[41]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85156.4]
  assign _T_509 = _GEN_3 >> _T_508; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85157.4]
  assign _T_511 = {io_a_data[42],io_data_in[42]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85159.4]
  assign _T_512 = _GEN_3 >> _T_511; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85160.4]
  assign _T_514 = {io_a_data[43],io_data_in[43]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85162.4]
  assign _T_515 = _GEN_3 >> _T_514; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85163.4]
  assign _T_517 = {io_a_data[44],io_data_in[44]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85165.4]
  assign _T_518 = _GEN_3 >> _T_517; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85166.4]
  assign _T_520 = {io_a_data[45],io_data_in[45]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85168.4]
  assign _T_521 = _GEN_3 >> _T_520; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85169.4]
  assign _T_523 = {io_a_data[46],io_data_in[46]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85171.4]
  assign _T_524 = _GEN_3 >> _T_523; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85172.4]
  assign _T_526 = {io_a_data[47],io_data_in[47]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85174.4]
  assign _T_527 = _GEN_3 >> _T_526; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85175.4]
  assign _T_529 = {io_a_data[48],io_data_in[48]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85177.4]
  assign _T_530 = _GEN_3 >> _T_529; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85178.4]
  assign _T_532 = {io_a_data[49],io_data_in[49]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85180.4]
  assign _T_533 = _GEN_3 >> _T_532; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85181.4]
  assign _T_535 = {io_a_data[50],io_data_in[50]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85183.4]
  assign _T_536 = _GEN_3 >> _T_535; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85184.4]
  assign _T_538 = {io_a_data[51],io_data_in[51]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85186.4]
  assign _T_539 = _GEN_3 >> _T_538; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85187.4]
  assign _T_541 = {io_a_data[52],io_data_in[52]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85189.4]
  assign _T_542 = _GEN_3 >> _T_541; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85190.4]
  assign _T_544 = {io_a_data[53],io_data_in[53]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85192.4]
  assign _T_545 = _GEN_3 >> _T_544; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85193.4]
  assign _T_547 = {io_a_data[54],io_data_in[54]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85195.4]
  assign _T_548 = _GEN_3 >> _T_547; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85196.4]
  assign _T_550 = {io_a_data[55],io_data_in[55]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85198.4]
  assign _T_551 = _GEN_3 >> _T_550; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85199.4]
  assign _T_553 = {io_a_data[56],io_data_in[56]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85201.4]
  assign _T_554 = _GEN_3 >> _T_553; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85202.4]
  assign _T_556 = {io_a_data[57],io_data_in[57]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85204.4]
  assign _T_557 = _GEN_3 >> _T_556; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85205.4]
  assign _T_559 = {io_a_data[58],io_data_in[58]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85207.4]
  assign _T_560 = _GEN_3 >> _T_559; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85208.4]
  assign _T_562 = {io_a_data[59],io_data_in[59]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85210.4]
  assign _T_563 = _GEN_3 >> _T_562; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85211.4]
  assign _T_565 = {io_a_data[60],io_data_in[60]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85213.4]
  assign _T_566 = _GEN_3 >> _T_565; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85214.4]
  assign _T_568 = {io_a_data[61],io_data_in[61]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85216.4]
  assign _T_569 = _GEN_3 >> _T_568; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85217.4]
  assign _T_571 = {io_a_data[62],io_data_in[62]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85219.4]
  assign _T_572 = _GEN_3 >> _T_571; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85220.4]
  assign _T_574 = {io_a_data[63],io_data_in[63]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85222.4]
  assign _T_575 = _GEN_3 >> _T_574; // @[Atomics.scala 44:8:chipyard.TestHarness.RocketConfig.fir@85223.4]
  assign _T_583 = {_T_407[0],_T_404[0],_T_401[0],_T_398[0],_T_395[0],_T_392[0],_T_389[0],_T_386[0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85231.4]
  assign _T_591 = {_T_431[0],_T_428[0],_T_425[0],_T_422[0],_T_419[0],_T_416[0],_T_413[0],_T_410[0],_T_583}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85239.4]
  assign _T_598 = {_T_455[0],_T_452[0],_T_449[0],_T_446[0],_T_443[0],_T_440[0],_T_437[0],_T_434[0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85246.4]
  assign _T_607 = {_T_479[0],_T_476[0],_T_473[0],_T_470[0],_T_467[0],_T_464[0],_T_461[0],_T_458[0],_T_598,_T_591}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85255.4]
  assign _T_614 = {_T_503[0],_T_500[0],_T_497[0],_T_494[0],_T_491[0],_T_488[0],_T_485[0],_T_482[0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85262.4]
  assign _T_622 = {_T_527[0],_T_524[0],_T_521[0],_T_518[0],_T_515[0],_T_512[0],_T_509[0],_T_506[0],_T_614}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85270.4]
  assign _T_629 = {_T_551[0],_T_548[0],_T_545[0],_T_542[0],_T_539[0],_T_536[0],_T_533[0],_T_530[0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85277.4]
  assign _T_638 = {_T_575[0],_T_572[0],_T_569[0],_T_566[0],_T_563[0],_T_560[0],_T_557[0],_T_554[0],_T_629,_T_622}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85286.4]
  assign logical = {_T_638,_T_607}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85287.4]
  assign _T_640 = adder ? 2'h2 : {{1'd0}, pick_a}; // @[Atomics.scala 51:8:chipyard.TestHarness.RocketConfig.fir@85289.4]
  assign _GEN_6 = 3'h2 == io_a_opcode ? _T_640 : 2'h1; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  assign _GEN_7 = 3'h3 == io_a_opcode ? 2'h3 : _GEN_6; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  assign _GEN_8 = 3'h4 == io_a_opcode ? 2'h0 : _GEN_7; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  assign _GEN_9 = 3'h5 == io_a_opcode ? 2'h0 : _GEN_8; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  assign _GEN_10 = 3'h6 == io_a_opcode ? 2'h0 : _GEN_9; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  assign _GEN_11 = 3'h7 == io_a_opcode ? 2'h0 : _GEN_10; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  assign select = io_write ? 2'h1 : _GEN_11; // @[Atomics.scala 48:19:chipyard.TestHarness.RocketConfig.fir@85300.4]
  assign selects_0 = io_a_mask[0] ? select : 2'h0; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85309.4]
  assign selects_1 = io_a_mask[1] ? select : 2'h0; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85310.4]
  assign selects_2 = io_a_mask[2] ? select : 2'h0; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85311.4]
  assign selects_3 = io_a_mask[3] ? select : 2'h0; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85312.4]
  assign selects_4 = io_a_mask[4] ? select : 2'h0; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85313.4]
  assign selects_5 = io_a_mask[5] ? select : 2'h0; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85314.4]
  assign selects_6 = io_a_mask[6] ? select : 2'h0; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85315.4]
  assign selects_7 = io_a_mask[7] ? select : 2'h0; // @[Atomics.scala 60:47:chipyard.TestHarness.RocketConfig.fir@85316.4]
  assign _GEN_13 = 2'h1 == selects_1 ? io_a_data[15:8] : io_data_in[15:8]; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85397.4]
  assign _GEN_14 = 2'h2 == selects_1 ? sum[15:8] : _GEN_13; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85397.4]
  assign _GEN_15 = 2'h3 == selects_1 ? logical[15:8] : _GEN_14; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85397.4]
  assign _GEN_17 = 2'h1 == selects_0 ? io_a_data[7:0] : io_data_in[7:0]; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85397.4]
  assign _GEN_18 = 2'h2 == selects_0 ? sum[7:0] : _GEN_17; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85397.4]
  assign _GEN_19 = 2'h3 == selects_0 ? logical[7:0] : _GEN_18; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85397.4]
  assign _GEN_21 = 2'h1 == selects_3 ? io_a_data[31:24] : io_data_in[31:24]; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85398.4]
  assign _GEN_22 = 2'h2 == selects_3 ? sum[31:24] : _GEN_21; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85398.4]
  assign _GEN_23 = 2'h3 == selects_3 ? logical[31:24] : _GEN_22; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85398.4]
  assign _GEN_25 = 2'h1 == selects_2 ? io_a_data[23:16] : io_data_in[23:16]; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85398.4]
  assign _GEN_26 = 2'h2 == selects_2 ? sum[23:16] : _GEN_25; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85398.4]
  assign _GEN_27 = 2'h3 == selects_2 ? logical[23:16] : _GEN_26; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85398.4]
  assign _T_692 = {_GEN_23,_GEN_27,_GEN_15,_GEN_19}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85399.4]
  assign _GEN_29 = 2'h1 == selects_5 ? io_a_data[47:40] : io_data_in[47:40]; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85400.4]
  assign _GEN_30 = 2'h2 == selects_5 ? sum[47:40] : _GEN_29; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85400.4]
  assign _GEN_31 = 2'h3 == selects_5 ? logical[47:40] : _GEN_30; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85400.4]
  assign _GEN_33 = 2'h1 == selects_4 ? io_a_data[39:32] : io_data_in[39:32]; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85400.4]
  assign _GEN_34 = 2'h2 == selects_4 ? sum[39:32] : _GEN_33; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85400.4]
  assign _GEN_35 = 2'h3 == selects_4 ? logical[39:32] : _GEN_34; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85400.4]
  assign _GEN_37 = 2'h1 == selects_7 ? io_a_data[63:56] : io_data_in[63:56]; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85401.4]
  assign _GEN_38 = 2'h2 == selects_7 ? sum[63:56] : _GEN_37; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85401.4]
  assign _GEN_39 = 2'h3 == selects_7 ? logical[63:56] : _GEN_38; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85401.4]
  assign _GEN_41 = 2'h1 == selects_6 ? io_a_data[55:48] : io_data_in[55:48]; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85401.4]
  assign _GEN_42 = 2'h2 == selects_6 ? sum[55:48] : _GEN_41; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85401.4]
  assign _GEN_43 = 2'h3 == selects_6 ? logical[55:48] : _GEN_42; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85401.4]
  assign _T_695 = {_GEN_39,_GEN_43,_GEN_31,_GEN_35}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@85402.4]
  assign io_data_out = {_T_695,_T_692}; // @[Atomics.scala 61:15:chipyard.TestHarness.RocketConfig.fir@85404.4]
endmodule
