module IntSyncCrossingSource( // @[:chipyard.TestHarness.RocketConfig.fir@129110.2]
  input   auto_in_0, // @[:chipyard.TestHarness.RocketConfig.fir@129113.4]
  output  auto_out_sync_0 // @[:chipyard.TestHarness.RocketConfig.fir@129113.4]
);
  assign auto_out_sync_0 = auto_in_0; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@129122.4]
endmodule
