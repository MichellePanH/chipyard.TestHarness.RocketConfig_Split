module IntXbar( // @[:chipyard.TestHarness.RocketConfig.fir@3.2]
  input   auto_int_in_0, // @[:chipyard.TestHarness.RocketConfig.fir@6.4]
  output  auto_int_out_0 // @[:chipyard.TestHarness.RocketConfig.fir@6.4]
);
  assign auto_int_out_0 = auto_int_in_0; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@15.4]
endmodule
