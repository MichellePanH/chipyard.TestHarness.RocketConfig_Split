module CompareRecFN( // @[:chipyard.TestHarness.RocketConfig.fir@234538.2]
  input  [64:0] io_a, // @[:chipyard.TestHarness.RocketConfig.fir@234539.4]
  input  [64:0] io_b, // @[:chipyard.TestHarness.RocketConfig.fir@234539.4]
  input         io_signaling, // @[:chipyard.TestHarness.RocketConfig.fir@234539.4]
  output        io_lt, // @[:chipyard.TestHarness.RocketConfig.fir@234539.4]
  output        io_eq, // @[:chipyard.TestHarness.RocketConfig.fir@234539.4]
  output [4:0]  io_exceptionFlags // @[:chipyard.TestHarness.RocketConfig.fir@234539.4]
);
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54:chipyard.TestHarness.RocketConfig.fir@234544.4]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54:chipyard.TestHarness.RocketConfig.fir@234546.4]
  wire  rawA_isNaN; // @[rawFloatFromRecFN.scala 55:33:chipyard.TestHarness.RocketConfig.fir@234550.4]
  wire  _T_8; // @[rawFloatFromRecFN.scala 56:36:chipyard.TestHarness.RocketConfig.fir@234553.4]
  wire  rawA_isInf; // @[rawFloatFromRecFN.scala 56:33:chipyard.TestHarness.RocketConfig.fir@234554.4]
  wire  rawA_sign; // @[rawFloatFromRecFN.scala 58:25:chipyard.TestHarness.RocketConfig.fir@234557.4]
  wire [12:0] rawA_sExp; // @[rawFloatFromRecFN.scala 59:27:chipyard.TestHarness.RocketConfig.fir@234559.4]
  wire  _T_12; // @[rawFloatFromRecFN.scala 60:39:chipyard.TestHarness.RocketConfig.fir@234561.4]
  wire [53:0] rawA_sig; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@234564.4]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54:chipyard.TestHarness.RocketConfig.fir@234568.4]
  wire  _T_20; // @[rawFloatFromRecFN.scala 52:54:chipyard.TestHarness.RocketConfig.fir@234570.4]
  wire  rawB_isNaN; // @[rawFloatFromRecFN.scala 55:33:chipyard.TestHarness.RocketConfig.fir@234574.4]
  wire  _T_24; // @[rawFloatFromRecFN.scala 56:36:chipyard.TestHarness.RocketConfig.fir@234577.4]
  wire  rawB_isInf; // @[rawFloatFromRecFN.scala 56:33:chipyard.TestHarness.RocketConfig.fir@234578.4]
  wire  rawB_sign; // @[rawFloatFromRecFN.scala 58:25:chipyard.TestHarness.RocketConfig.fir@234581.4]
  wire [12:0] rawB_sExp; // @[rawFloatFromRecFN.scala 59:27:chipyard.TestHarness.RocketConfig.fir@234583.4]
  wire  _T_28; // @[rawFloatFromRecFN.scala 60:39:chipyard.TestHarness.RocketConfig.fir@234585.4]
  wire [53:0] rawB_sig; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@234588.4]
  wire  _T_32; // @[CompareRecFN.scala 57:19:chipyard.TestHarness.RocketConfig.fir@234590.4]
  wire  _T_33; // @[CompareRecFN.scala 57:35:chipyard.TestHarness.RocketConfig.fir@234591.4]
  wire  ordered; // @[CompareRecFN.scala 57:32:chipyard.TestHarness.RocketConfig.fir@234592.4]
  wire  bothInfs; // @[CompareRecFN.scala 58:33:chipyard.TestHarness.RocketConfig.fir@234593.4]
  wire  bothZeros; // @[CompareRecFN.scala 59:33:chipyard.TestHarness.RocketConfig.fir@234594.4]
  wire  eqExps; // @[CompareRecFN.scala 60:29:chipyard.TestHarness.RocketConfig.fir@234595.4]
  wire  _T_34; // @[CompareRecFN.scala 62:20:chipyard.TestHarness.RocketConfig.fir@234596.4]
  wire  _T_35; // @[CompareRecFN.scala 62:57:chipyard.TestHarness.RocketConfig.fir@234597.4]
  wire  _T_36; // @[CompareRecFN.scala 62:44:chipyard.TestHarness.RocketConfig.fir@234598.4]
  wire  common_ltMags; // @[CompareRecFN.scala 62:33:chipyard.TestHarness.RocketConfig.fir@234599.4]
  wire  _T_37; // @[CompareRecFN.scala 63:45:chipyard.TestHarness.RocketConfig.fir@234600.4]
  wire  common_eqMags; // @[CompareRecFN.scala 63:32:chipyard.TestHarness.RocketConfig.fir@234601.4]
  wire  _T_38; // @[CompareRecFN.scala 66:9:chipyard.TestHarness.RocketConfig.fir@234602.4]
  wire  _T_39; // @[CompareRecFN.scala 67:28:chipyard.TestHarness.RocketConfig.fir@234603.4]
  wire  _T_40; // @[CompareRecFN.scala 67:25:chipyard.TestHarness.RocketConfig.fir@234604.4]
  wire  _T_41; // @[CompareRecFN.scala 68:19:chipyard.TestHarness.RocketConfig.fir@234605.4]
  wire  _T_42; // @[CompareRecFN.scala 69:38:chipyard.TestHarness.RocketConfig.fir@234606.4]
  wire  _T_43; // @[CompareRecFN.scala 69:35:chipyard.TestHarness.RocketConfig.fir@234607.4]
  wire  _T_44; // @[CompareRecFN.scala 69:57:chipyard.TestHarness.RocketConfig.fir@234608.4]
  wire  _T_45; // @[CompareRecFN.scala 69:54:chipyard.TestHarness.RocketConfig.fir@234609.4]
  wire  _T_47; // @[CompareRecFN.scala 70:41:chipyard.TestHarness.RocketConfig.fir@234611.4]
  wire  _T_48; // @[CompareRecFN.scala 69:74:chipyard.TestHarness.RocketConfig.fir@234612.4]
  wire  _T_49; // @[CompareRecFN.scala 68:30:chipyard.TestHarness.RocketConfig.fir@234613.4]
  wire  _T_50; // @[CompareRecFN.scala 67:41:chipyard.TestHarness.RocketConfig.fir@234614.4]
  wire  ordered_lt; // @[CompareRecFN.scala 66:21:chipyard.TestHarness.RocketConfig.fir@234615.4]
  wire  _T_51; // @[CompareRecFN.scala 72:34:chipyard.TestHarness.RocketConfig.fir@234616.4]
  wire  _T_52; // @[CompareRecFN.scala 72:62:chipyard.TestHarness.RocketConfig.fir@234617.4]
  wire  _T_53; // @[CompareRecFN.scala 72:49:chipyard.TestHarness.RocketConfig.fir@234618.4]
  wire  ordered_eq; // @[CompareRecFN.scala 72:19:chipyard.TestHarness.RocketConfig.fir@234619.4]
  wire  _T_55; // @[common.scala 81:49:chipyard.TestHarness.RocketConfig.fir@234621.4]
  wire  _T_56; // @[common.scala 81:46:chipyard.TestHarness.RocketConfig.fir@234622.4]
  wire  _T_58; // @[common.scala 81:49:chipyard.TestHarness.RocketConfig.fir@234624.4]
  wire  _T_59; // @[common.scala 81:46:chipyard.TestHarness.RocketConfig.fir@234625.4]
  wire  _T_60; // @[CompareRecFN.scala 75:32:chipyard.TestHarness.RocketConfig.fir@234626.4]
  wire  _T_61; // @[CompareRecFN.scala 76:30:chipyard.TestHarness.RocketConfig.fir@234627.4]
  wire  _T_62; // @[CompareRecFN.scala 76:27:chipyard.TestHarness.RocketConfig.fir@234628.4]
  wire  invalid; // @[CompareRecFN.scala 75:58:chipyard.TestHarness.RocketConfig.fir@234629.4]
  assign rawA_isZero = io_a[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54:chipyard.TestHarness.RocketConfig.fir@234544.4]
  assign _T_4 = io_a[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54:chipyard.TestHarness.RocketConfig.fir@234546.4]
  assign rawA_isNaN = _T_4 & io_a[61]; // @[rawFloatFromRecFN.scala 55:33:chipyard.TestHarness.RocketConfig.fir@234550.4]
  assign _T_8 = ~io_a[61]; // @[rawFloatFromRecFN.scala 56:36:chipyard.TestHarness.RocketConfig.fir@234553.4]
  assign rawA_isInf = _T_4 & _T_8; // @[rawFloatFromRecFN.scala 56:33:chipyard.TestHarness.RocketConfig.fir@234554.4]
  assign rawA_sign = io_a[64]; // @[rawFloatFromRecFN.scala 58:25:chipyard.TestHarness.RocketConfig.fir@234557.4]
  assign rawA_sExp = {1'b0,$signed(io_a[63:52])}; // @[rawFloatFromRecFN.scala 59:27:chipyard.TestHarness.RocketConfig.fir@234559.4]
  assign _T_12 = ~rawA_isZero; // @[rawFloatFromRecFN.scala 60:39:chipyard.TestHarness.RocketConfig.fir@234561.4]
  assign rawA_sig = {1'h0,_T_12,io_a[51:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@234564.4]
  assign rawB_isZero = io_b[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54:chipyard.TestHarness.RocketConfig.fir@234568.4]
  assign _T_20 = io_b[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54:chipyard.TestHarness.RocketConfig.fir@234570.4]
  assign rawB_isNaN = _T_20 & io_b[61]; // @[rawFloatFromRecFN.scala 55:33:chipyard.TestHarness.RocketConfig.fir@234574.4]
  assign _T_24 = ~io_b[61]; // @[rawFloatFromRecFN.scala 56:36:chipyard.TestHarness.RocketConfig.fir@234577.4]
  assign rawB_isInf = _T_20 & _T_24; // @[rawFloatFromRecFN.scala 56:33:chipyard.TestHarness.RocketConfig.fir@234578.4]
  assign rawB_sign = io_b[64]; // @[rawFloatFromRecFN.scala 58:25:chipyard.TestHarness.RocketConfig.fir@234581.4]
  assign rawB_sExp = {1'b0,$signed(io_b[63:52])}; // @[rawFloatFromRecFN.scala 59:27:chipyard.TestHarness.RocketConfig.fir@234583.4]
  assign _T_28 = ~rawB_isZero; // @[rawFloatFromRecFN.scala 60:39:chipyard.TestHarness.RocketConfig.fir@234585.4]
  assign rawB_sig = {1'h0,_T_28,io_b[51:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@234588.4]
  assign _T_32 = ~rawA_isNaN; // @[CompareRecFN.scala 57:19:chipyard.TestHarness.RocketConfig.fir@234590.4]
  assign _T_33 = ~rawB_isNaN; // @[CompareRecFN.scala 57:35:chipyard.TestHarness.RocketConfig.fir@234591.4]
  assign ordered = _T_32 & _T_33; // @[CompareRecFN.scala 57:32:chipyard.TestHarness.RocketConfig.fir@234592.4]
  assign bothInfs = rawA_isInf & rawB_isInf; // @[CompareRecFN.scala 58:33:chipyard.TestHarness.RocketConfig.fir@234593.4]
  assign bothZeros = rawA_isZero & rawB_isZero; // @[CompareRecFN.scala 59:33:chipyard.TestHarness.RocketConfig.fir@234594.4]
  assign eqExps = $signed(rawA_sExp) == $signed(rawB_sExp); // @[CompareRecFN.scala 60:29:chipyard.TestHarness.RocketConfig.fir@234595.4]
  assign _T_34 = $signed(rawA_sExp) < $signed(rawB_sExp); // @[CompareRecFN.scala 62:20:chipyard.TestHarness.RocketConfig.fir@234596.4]
  assign _T_35 = rawA_sig < rawB_sig; // @[CompareRecFN.scala 62:57:chipyard.TestHarness.RocketConfig.fir@234597.4]
  assign _T_36 = eqExps & _T_35; // @[CompareRecFN.scala 62:44:chipyard.TestHarness.RocketConfig.fir@234598.4]
  assign common_ltMags = _T_34 | _T_36; // @[CompareRecFN.scala 62:33:chipyard.TestHarness.RocketConfig.fir@234599.4]
  assign _T_37 = rawA_sig == rawB_sig; // @[CompareRecFN.scala 63:45:chipyard.TestHarness.RocketConfig.fir@234600.4]
  assign common_eqMags = eqExps & _T_37; // @[CompareRecFN.scala 63:32:chipyard.TestHarness.RocketConfig.fir@234601.4]
  assign _T_38 = ~bothZeros; // @[CompareRecFN.scala 66:9:chipyard.TestHarness.RocketConfig.fir@234602.4]
  assign _T_39 = ~rawB_sign; // @[CompareRecFN.scala 67:28:chipyard.TestHarness.RocketConfig.fir@234603.4]
  assign _T_40 = rawA_sign & _T_39; // @[CompareRecFN.scala 67:25:chipyard.TestHarness.RocketConfig.fir@234604.4]
  assign _T_41 = ~bothInfs; // @[CompareRecFN.scala 68:19:chipyard.TestHarness.RocketConfig.fir@234605.4]
  assign _T_42 = ~common_ltMags; // @[CompareRecFN.scala 69:38:chipyard.TestHarness.RocketConfig.fir@234606.4]
  assign _T_43 = rawA_sign & _T_42; // @[CompareRecFN.scala 69:35:chipyard.TestHarness.RocketConfig.fir@234607.4]
  assign _T_44 = ~common_eqMags; // @[CompareRecFN.scala 69:57:chipyard.TestHarness.RocketConfig.fir@234608.4]
  assign _T_45 = _T_43 & _T_44; // @[CompareRecFN.scala 69:54:chipyard.TestHarness.RocketConfig.fir@234609.4]
  assign _T_47 = _T_39 & common_ltMags; // @[CompareRecFN.scala 70:41:chipyard.TestHarness.RocketConfig.fir@234611.4]
  assign _T_48 = _T_45 | _T_47; // @[CompareRecFN.scala 69:74:chipyard.TestHarness.RocketConfig.fir@234612.4]
  assign _T_49 = _T_41 & _T_48; // @[CompareRecFN.scala 68:30:chipyard.TestHarness.RocketConfig.fir@234613.4]
  assign _T_50 = _T_40 | _T_49; // @[CompareRecFN.scala 67:41:chipyard.TestHarness.RocketConfig.fir@234614.4]
  assign ordered_lt = _T_38 & _T_50; // @[CompareRecFN.scala 66:21:chipyard.TestHarness.RocketConfig.fir@234615.4]
  assign _T_51 = rawA_sign == rawB_sign; // @[CompareRecFN.scala 72:34:chipyard.TestHarness.RocketConfig.fir@234616.4]
  assign _T_52 = bothInfs | common_eqMags; // @[CompareRecFN.scala 72:62:chipyard.TestHarness.RocketConfig.fir@234617.4]
  assign _T_53 = _T_51 & _T_52; // @[CompareRecFN.scala 72:49:chipyard.TestHarness.RocketConfig.fir@234618.4]
  assign ordered_eq = bothZeros | _T_53; // @[CompareRecFN.scala 72:19:chipyard.TestHarness.RocketConfig.fir@234619.4]
  assign _T_55 = ~rawA_sig[51]; // @[common.scala 81:49:chipyard.TestHarness.RocketConfig.fir@234621.4]
  assign _T_56 = rawA_isNaN & _T_55; // @[common.scala 81:46:chipyard.TestHarness.RocketConfig.fir@234622.4]
  assign _T_58 = ~rawB_sig[51]; // @[common.scala 81:49:chipyard.TestHarness.RocketConfig.fir@234624.4]
  assign _T_59 = rawB_isNaN & _T_58; // @[common.scala 81:46:chipyard.TestHarness.RocketConfig.fir@234625.4]
  assign _T_60 = _T_56 | _T_59; // @[CompareRecFN.scala 75:32:chipyard.TestHarness.RocketConfig.fir@234626.4]
  assign _T_61 = ~ordered; // @[CompareRecFN.scala 76:30:chipyard.TestHarness.RocketConfig.fir@234627.4]
  assign _T_62 = io_signaling & _T_61; // @[CompareRecFN.scala 76:27:chipyard.TestHarness.RocketConfig.fir@234628.4]
  assign invalid = _T_60 | _T_62; // @[CompareRecFN.scala 75:58:chipyard.TestHarness.RocketConfig.fir@234629.4]
  assign io_lt = ordered & ordered_lt; // @[CompareRecFN.scala 78:11:chipyard.TestHarness.RocketConfig.fir@234631.4]
  assign io_eq = ordered & ordered_eq; // @[CompareRecFN.scala 79:11:chipyard.TestHarness.RocketConfig.fir@234633.4]
  assign io_exceptionFlags = {invalid,4'h0}; // @[CompareRecFN.scala 81:23:chipyard.TestHarness.RocketConfig.fir@234640.4]
endmodule
