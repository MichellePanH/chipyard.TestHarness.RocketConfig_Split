module TLFIFOFixer( // @[:chipyard.TestHarness.RocketConfig.fir@10931.2]
  input         clock, // @[:chipyard.TestHarness.RocketConfig.fir@10932.4]
  input         reset, // @[:chipyard.TestHarness.RocketConfig.fir@10933.4]
  output        auto_in_1_a_ready, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_in_1_a_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [2:0]  auto_in_1_a_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [2:0]  auto_in_1_a_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [3:0]  auto_in_1_a_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [1:0]  auto_in_1_a_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [31:0] auto_in_1_a_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [7:0]  auto_in_1_a_bits_mask, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [63:0] auto_in_1_a_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_in_1_a_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_in_1_b_ready, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_in_1_b_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [1:0]  auto_in_1_b_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [31:0] auto_in_1_b_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_in_1_c_ready, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_in_1_c_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [2:0]  auto_in_1_c_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [2:0]  auto_in_1_c_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [3:0]  auto_in_1_c_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [1:0]  auto_in_1_c_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [31:0] auto_in_1_c_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [63:0] auto_in_1_c_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_in_1_c_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_in_1_d_ready, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_in_1_d_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [2:0]  auto_in_1_d_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [1:0]  auto_in_1_d_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [3:0]  auto_in_1_d_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [1:0]  auto_in_1_d_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [2:0]  auto_in_1_d_bits_sink, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_in_1_d_bits_denied, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [63:0] auto_in_1_d_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_in_1_d_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_in_1_e_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [2:0]  auto_in_1_e_bits_sink, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_in_0_a_ready, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_in_0_a_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [2:0]  auto_in_0_a_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [2:0]  auto_in_0_a_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [3:0]  auto_in_0_a_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_in_0_a_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [31:0] auto_in_0_a_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [7:0]  auto_in_0_a_bits_mask, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [63:0] auto_in_0_a_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_in_0_a_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_in_0_d_ready, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_in_0_d_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [2:0]  auto_in_0_d_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [1:0]  auto_in_0_d_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [3:0]  auto_in_0_d_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [2:0]  auto_in_0_d_bits_sink, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_in_0_d_bits_denied, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [63:0] auto_in_0_d_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_in_0_d_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_out_1_a_ready, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_out_1_a_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [2:0]  auto_out_1_a_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [2:0]  auto_out_1_a_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [3:0]  auto_out_1_a_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [1:0]  auto_out_1_a_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [31:0] auto_out_1_a_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [7:0]  auto_out_1_a_bits_mask, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [63:0] auto_out_1_a_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_out_1_a_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_out_1_b_ready, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_out_1_b_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [1:0]  auto_out_1_b_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [31:0] auto_out_1_b_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_out_1_c_ready, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_out_1_c_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [2:0]  auto_out_1_c_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [2:0]  auto_out_1_c_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [3:0]  auto_out_1_c_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [1:0]  auto_out_1_c_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [31:0] auto_out_1_c_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [63:0] auto_out_1_c_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_out_1_c_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_out_1_d_ready, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_out_1_d_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [2:0]  auto_out_1_d_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [1:0]  auto_out_1_d_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [3:0]  auto_out_1_d_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [1:0]  auto_out_1_d_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [2:0]  auto_out_1_d_bits_sink, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_out_1_d_bits_denied, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [63:0] auto_out_1_d_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_out_1_d_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_out_1_e_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [2:0]  auto_out_1_e_bits_sink, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_out_0_a_ready, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_out_0_a_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [2:0]  auto_out_0_a_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [2:0]  auto_out_0_a_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [3:0]  auto_out_0_a_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_out_0_a_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [31:0] auto_out_0_a_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [7:0]  auto_out_0_a_bits_mask, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output [63:0] auto_out_0_a_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_out_0_a_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  output        auto_out_0_d_ready, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_out_0_d_valid, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [2:0]  auto_out_0_d_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [1:0]  auto_out_0_d_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [3:0]  auto_out_0_d_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [2:0]  auto_out_0_d_bits_sink, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_out_0_d_bits_denied, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input  [63:0] auto_out_0_d_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
  input         auto_out_0_d_bits_corrupt // @[:chipyard.TestHarness.RocketConfig.fir@10934.4]
);
  wire  TLMonitor_clock; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire  TLMonitor_reset; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire  TLMonitor_io_in_a_ready; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire  TLMonitor_io_in_a_valid; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire [2:0] TLMonitor_io_in_a_bits_opcode; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire [2:0] TLMonitor_io_in_a_bits_param; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire [3:0] TLMonitor_io_in_a_bits_size; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire  TLMonitor_io_in_a_bits_source; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire [31:0] TLMonitor_io_in_a_bits_address; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire [7:0] TLMonitor_io_in_a_bits_mask; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire  TLMonitor_io_in_a_bits_corrupt; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire  TLMonitor_io_in_d_ready; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire  TLMonitor_io_in_d_valid; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire [2:0] TLMonitor_io_in_d_bits_opcode; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire [1:0] TLMonitor_io_in_d_bits_param; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire [3:0] TLMonitor_io_in_d_bits_size; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire [2:0] TLMonitor_io_in_d_bits_sink; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire  TLMonitor_io_in_d_bits_denied; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire  TLMonitor_io_in_d_bits_corrupt; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
  wire  TLMonitor_1_clock; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_reset; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_io_in_a_ready; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_io_in_a_valid; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [2:0] TLMonitor_1_io_in_a_bits_opcode; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [2:0] TLMonitor_1_io_in_a_bits_param; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [3:0] TLMonitor_1_io_in_a_bits_size; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [1:0] TLMonitor_1_io_in_a_bits_source; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [31:0] TLMonitor_1_io_in_a_bits_address; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [7:0] TLMonitor_1_io_in_a_bits_mask; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_io_in_a_bits_corrupt; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_io_in_b_ready; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_io_in_b_valid; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [1:0] TLMonitor_1_io_in_b_bits_param; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [31:0] TLMonitor_1_io_in_b_bits_address; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_io_in_c_ready; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_io_in_c_valid; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [2:0] TLMonitor_1_io_in_c_bits_opcode; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [2:0] TLMonitor_1_io_in_c_bits_param; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [3:0] TLMonitor_1_io_in_c_bits_size; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [1:0] TLMonitor_1_io_in_c_bits_source; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [31:0] TLMonitor_1_io_in_c_bits_address; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_io_in_c_bits_corrupt; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_io_in_d_ready; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_io_in_d_valid; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [2:0] TLMonitor_1_io_in_d_bits_opcode; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [1:0] TLMonitor_1_io_in_d_bits_param; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [3:0] TLMonitor_1_io_in_d_bits_size; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [1:0] TLMonitor_1_io_in_d_bits_source; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [2:0] TLMonitor_1_io_in_d_bits_sink; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_io_in_d_bits_denied; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_io_in_d_bits_corrupt; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire  TLMonitor_1_io_in_e_valid; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  wire [2:0] TLMonitor_1_io_in_e_bits_sink; // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
  TLMonitor_2 TLMonitor ( // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10943.4]
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt)
  );
  TLMonitor_3 TLMonitor_1 ( // @[Nodes.scala 25:25:chipyard.TestHarness.RocketConfig.fir@10966.4]
    .clock(TLMonitor_1_clock),
    .reset(TLMonitor_1_reset),
    .io_in_a_ready(TLMonitor_1_io_in_a_ready),
    .io_in_a_valid(TLMonitor_1_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_1_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_1_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_1_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_1_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_1_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_1_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_1_io_in_a_bits_corrupt),
    .io_in_b_ready(TLMonitor_1_io_in_b_ready),
    .io_in_b_valid(TLMonitor_1_io_in_b_valid),
    .io_in_b_bits_param(TLMonitor_1_io_in_b_bits_param),
    .io_in_b_bits_address(TLMonitor_1_io_in_b_bits_address),
    .io_in_c_ready(TLMonitor_1_io_in_c_ready),
    .io_in_c_valid(TLMonitor_1_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_1_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_1_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_1_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_1_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_1_io_in_c_bits_address),
    .io_in_c_bits_corrupt(TLMonitor_1_io_in_c_bits_corrupt),
    .io_in_d_ready(TLMonitor_1_io_in_d_ready),
    .io_in_d_valid(TLMonitor_1_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_1_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_1_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_1_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_1_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_1_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_1_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_1_io_in_d_bits_corrupt),
    .io_in_e_valid(TLMonitor_1_io_in_e_valid),
    .io_in_e_bits_sink(TLMonitor_1_io_in_e_bits_sink)
  );
  assign auto_in_1_a_ready = auto_out_1_a_ready; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_1_b_valid = auto_out_1_b_valid; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_1_b_bits_param = auto_out_1_b_bits_param; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_1_b_bits_address = auto_out_1_b_bits_address; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_1_c_ready = auto_out_1_c_ready; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_1_d_valid = auto_out_1_d_valid; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_1_d_bits_opcode = auto_out_1_d_bits_opcode; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_1_d_bits_param = auto_out_1_d_bits_param; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_1_d_bits_size = auto_out_1_d_bits_size; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_1_d_bits_source = auto_out_1_d_bits_source; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_1_d_bits_sink = auto_out_1_d_bits_sink; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_1_d_bits_denied = auto_out_1_d_bits_denied; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_1_d_bits_data = auto_out_1_d_bits_data; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_1_d_bits_corrupt = auto_out_1_d_bits_corrupt; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11018.4]
  assign auto_in_0_a_ready = auto_out_0_a_ready; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11017.4]
  assign auto_in_0_d_valid = auto_out_0_d_valid; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11017.4]
  assign auto_in_0_d_bits_opcode = auto_out_0_d_bits_opcode; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11017.4]
  assign auto_in_0_d_bits_param = auto_out_0_d_bits_param; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11017.4]
  assign auto_in_0_d_bits_size = auto_out_0_d_bits_size; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11017.4]
  assign auto_in_0_d_bits_sink = auto_out_0_d_bits_sink; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11017.4]
  assign auto_in_0_d_bits_denied = auto_out_0_d_bits_denied; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11017.4]
  assign auto_in_0_d_bits_data = auto_out_0_d_bits_data; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11017.4]
  assign auto_in_0_d_bits_corrupt = auto_out_0_d_bits_corrupt; // @[LazyModule.scala 181:31:chipyard.TestHarness.RocketConfig.fir@11017.4]
  assign auto_out_1_a_valid = auto_in_1_a_valid; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_a_bits_opcode = auto_in_1_a_bits_opcode; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_a_bits_param = auto_in_1_a_bits_param; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_a_bits_size = auto_in_1_a_bits_size; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_a_bits_source = auto_in_1_a_bits_source; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_a_bits_address = auto_in_1_a_bits_address; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_a_bits_mask = auto_in_1_a_bits_mask; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_a_bits_data = auto_in_1_a_bits_data; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_a_bits_corrupt = auto_in_1_a_bits_corrupt; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_b_ready = auto_in_1_b_ready; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_c_valid = auto_in_1_c_valid; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_c_bits_opcode = auto_in_1_c_bits_opcode; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_c_bits_param = auto_in_1_c_bits_param; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_c_bits_size = auto_in_1_c_bits_size; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_c_bits_source = auto_in_1_c_bits_source; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_c_bits_address = auto_in_1_c_bits_address; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_c_bits_data = auto_in_1_c_bits_data; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_c_bits_corrupt = auto_in_1_c_bits_corrupt; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_d_ready = auto_in_1_d_ready; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_e_valid = auto_in_1_e_valid; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_1_e_bits_sink = auto_in_1_e_bits_sink; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11016.4]
  assign auto_out_0_a_valid = auto_in_0_a_valid; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11015.4]
  assign auto_out_0_a_bits_opcode = auto_in_0_a_bits_opcode; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11015.4]
  assign auto_out_0_a_bits_param = auto_in_0_a_bits_param; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11015.4]
  assign auto_out_0_a_bits_size = auto_in_0_a_bits_size; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11015.4]
  assign auto_out_0_a_bits_source = auto_in_0_a_bits_source; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11015.4]
  assign auto_out_0_a_bits_address = auto_in_0_a_bits_address; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11015.4]
  assign auto_out_0_a_bits_mask = auto_in_0_a_bits_mask; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11015.4]
  assign auto_out_0_a_bits_data = auto_in_0_a_bits_data; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11015.4]
  assign auto_out_0_a_bits_corrupt = auto_in_0_a_bits_corrupt; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11015.4]
  assign auto_out_0_d_ready = auto_in_0_d_ready; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@11015.4]
  assign TLMonitor_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@10944.4]
  assign TLMonitor_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@10945.4]
  assign TLMonitor_io_in_a_ready = auto_out_0_a_ready; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10965.4]
  assign TLMonitor_io_in_a_valid = auto_in_0_a_valid; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10964.4]
  assign TLMonitor_io_in_a_bits_opcode = auto_in_0_a_bits_opcode; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10963.4]
  assign TLMonitor_io_in_a_bits_param = auto_in_0_a_bits_param; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10962.4]
  assign TLMonitor_io_in_a_bits_size = auto_in_0_a_bits_size; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10961.4]
  assign TLMonitor_io_in_a_bits_source = auto_in_0_a_bits_source; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10960.4]
  assign TLMonitor_io_in_a_bits_address = auto_in_0_a_bits_address; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10959.4]
  assign TLMonitor_io_in_a_bits_mask = auto_in_0_a_bits_mask; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10958.4]
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_0_a_bits_corrupt; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10956.4]
  assign TLMonitor_io_in_d_ready = auto_in_0_d_ready; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10955.4]
  assign TLMonitor_io_in_d_valid = auto_out_0_d_valid; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10954.4]
  assign TLMonitor_io_in_d_bits_opcode = auto_out_0_d_bits_opcode; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10953.4]
  assign TLMonitor_io_in_d_bits_param = auto_out_0_d_bits_param; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10952.4]
  assign TLMonitor_io_in_d_bits_size = auto_out_0_d_bits_size; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10951.4]
  assign TLMonitor_io_in_d_bits_sink = auto_out_0_d_bits_sink; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10949.4]
  assign TLMonitor_io_in_d_bits_denied = auto_out_0_d_bits_denied; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10948.4]
  assign TLMonitor_io_in_d_bits_corrupt = auto_out_0_d_bits_corrupt; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10946.4]
  assign TLMonitor_1_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@10967.4]
  assign TLMonitor_1_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@10968.4]
  assign TLMonitor_1_io_in_a_ready = auto_out_1_a_ready; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@11010.4]
  assign TLMonitor_1_io_in_a_valid = auto_in_1_a_valid; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@11009.4]
  assign TLMonitor_1_io_in_a_bits_opcode = auto_in_1_a_bits_opcode; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@11008.4]
  assign TLMonitor_1_io_in_a_bits_param = auto_in_1_a_bits_param; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@11007.4]
  assign TLMonitor_1_io_in_a_bits_size = auto_in_1_a_bits_size; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@11006.4]
  assign TLMonitor_1_io_in_a_bits_source = auto_in_1_a_bits_source; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@11005.4]
  assign TLMonitor_1_io_in_a_bits_address = auto_in_1_a_bits_address; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@11004.4]
  assign TLMonitor_1_io_in_a_bits_mask = auto_in_1_a_bits_mask; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@11003.4]
  assign TLMonitor_1_io_in_a_bits_corrupt = auto_in_1_a_bits_corrupt; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@11001.4]
  assign TLMonitor_1_io_in_b_ready = auto_in_1_b_ready; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@11000.4]
  assign TLMonitor_1_io_in_b_valid = auto_out_1_b_valid; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10999.4]
  assign TLMonitor_1_io_in_b_bits_param = auto_out_1_b_bits_param; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10997.4]
  assign TLMonitor_1_io_in_b_bits_address = auto_out_1_b_bits_address; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10994.4]
  assign TLMonitor_1_io_in_c_ready = auto_out_1_c_ready; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10990.4]
  assign TLMonitor_1_io_in_c_valid = auto_in_1_c_valid; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10989.4]
  assign TLMonitor_1_io_in_c_bits_opcode = auto_in_1_c_bits_opcode; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10988.4]
  assign TLMonitor_1_io_in_c_bits_param = auto_in_1_c_bits_param; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10987.4]
  assign TLMonitor_1_io_in_c_bits_size = auto_in_1_c_bits_size; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10986.4]
  assign TLMonitor_1_io_in_c_bits_source = auto_in_1_c_bits_source; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10985.4]
  assign TLMonitor_1_io_in_c_bits_address = auto_in_1_c_bits_address; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10984.4]
  assign TLMonitor_1_io_in_c_bits_corrupt = auto_in_1_c_bits_corrupt; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10982.4]
  assign TLMonitor_1_io_in_d_ready = auto_in_1_d_ready; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10981.4]
  assign TLMonitor_1_io_in_d_valid = auto_out_1_d_valid; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10980.4]
  assign TLMonitor_1_io_in_d_bits_opcode = auto_out_1_d_bits_opcode; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10979.4]
  assign TLMonitor_1_io_in_d_bits_param = auto_out_1_d_bits_param; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10978.4]
  assign TLMonitor_1_io_in_d_bits_size = auto_out_1_d_bits_size; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10977.4]
  assign TLMonitor_1_io_in_d_bits_source = auto_out_1_d_bits_source; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10976.4]
  assign TLMonitor_1_io_in_d_bits_sink = auto_out_1_d_bits_sink; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10975.4]
  assign TLMonitor_1_io_in_d_bits_denied = auto_out_1_d_bits_denied; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10974.4]
  assign TLMonitor_1_io_in_d_bits_corrupt = auto_out_1_d_bits_corrupt; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10972.4]
  assign TLMonitor_1_io_in_e_valid = auto_in_1_e_valid; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10970.4]
  assign TLMonitor_1_io_in_e_bits_sink = auto_in_1_e_bits_sink; // @[Nodes.scala 26:19:chipyard.TestHarness.RocketConfig.fir@10969.4]
endmodule
