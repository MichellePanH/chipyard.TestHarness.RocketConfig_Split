module BreakpointUnit( // @[:chipyard.TestHarness.RocketConfig.fir@249410.2]
  input         io_status_debug, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  input  [1:0]  io_status_prv, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  input         io_bp_0_control_action, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  input  [1:0]  io_bp_0_control_tmatch, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  input         io_bp_0_control_m, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  input         io_bp_0_control_s, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  input         io_bp_0_control_u, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  input         io_bp_0_control_x, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  input         io_bp_0_control_w, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  input         io_bp_0_control_r, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  input  [38:0] io_bp_0_address, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  input  [38:0] io_pc, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  input  [38:0] io_ea, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  output        io_xcpt_if, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  output        io_xcpt_ld, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  output        io_xcpt_st, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  output        io_debug_if, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  output        io_debug_ld, // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
  output        io_debug_st // @[:chipyard.TestHarness.RocketConfig.fir@249413.4]
);
  wire  _T; // @[Breakpoint.scala 31:35:chipyard.TestHarness.RocketConfig.fir@249421.4]
  wire [3:0] _T_3; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@249424.4]
  wire [3:0] _T_4; // @[Breakpoint.scala 31:68:chipyard.TestHarness.RocketConfig.fir@249425.4]
  wire  _T_6; // @[Breakpoint.scala 31:50:chipyard.TestHarness.RocketConfig.fir@249427.4]
  wire  _T_7; // @[Breakpoint.scala 83:16:chipyard.TestHarness.RocketConfig.fir@249428.4]
  wire  _T_9; // @[Breakpoint.scala 45:8:chipyard.TestHarness.RocketConfig.fir@249430.4]
  wire  _T_11; // @[Breakpoint.scala 45:20:chipyard.TestHarness.RocketConfig.fir@249432.4]
  wire [38:0] _T_12; // @[Breakpoint.scala 42:6:chipyard.TestHarness.RocketConfig.fir@249433.4]
  wire  _T_15; // @[Breakpoint.scala 39:73:chipyard.TestHarness.RocketConfig.fir@249436.4]
  wire  _T_17; // @[Breakpoint.scala 39:73:chipyard.TestHarness.RocketConfig.fir@249438.4]
  wire  _T_19; // @[Breakpoint.scala 39:73:chipyard.TestHarness.RocketConfig.fir@249440.4]
  wire [3:0] _T_22; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@249443.4]
  wire [38:0] _GEN_11; // @[Breakpoint.scala 42:9:chipyard.TestHarness.RocketConfig.fir@249444.4]
  wire [38:0] _T_23; // @[Breakpoint.scala 42:9:chipyard.TestHarness.RocketConfig.fir@249444.4]
  wire [38:0] _T_24; // @[Breakpoint.scala 42:24:chipyard.TestHarness.RocketConfig.fir@249445.4]
  wire [38:0] _T_35; // @[Breakpoint.scala 42:33:chipyard.TestHarness.RocketConfig.fir@249456.4]
  wire  _T_36; // @[Breakpoint.scala 42:19:chipyard.TestHarness.RocketConfig.fir@249457.4]
  wire  _T_37; // @[Breakpoint.scala 48:8:chipyard.TestHarness.RocketConfig.fir@249458.4]
  wire  _T_38; // @[Breakpoint.scala 83:32:chipyard.TestHarness.RocketConfig.fir@249459.4]
  wire  _T_39; // @[Breakpoint.scala 84:16:chipyard.TestHarness.RocketConfig.fir@249460.4]
  wire  _T_70; // @[Breakpoint.scala 84:32:chipyard.TestHarness.RocketConfig.fir@249491.4]
  wire  _T_71; // @[Breakpoint.scala 85:16:chipyard.TestHarness.RocketConfig.fir@249492.4]
  wire  _T_73; // @[Breakpoint.scala 45:8:chipyard.TestHarness.RocketConfig.fir@249494.4]
  wire  _T_75; // @[Breakpoint.scala 45:20:chipyard.TestHarness.RocketConfig.fir@249496.4]
  wire [38:0] _T_76; // @[Breakpoint.scala 42:6:chipyard.TestHarness.RocketConfig.fir@249497.4]
  wire [38:0] _T_87; // @[Breakpoint.scala 42:9:chipyard.TestHarness.RocketConfig.fir@249508.4]
  wire  _T_100; // @[Breakpoint.scala 42:19:chipyard.TestHarness.RocketConfig.fir@249521.4]
  wire  _T_101; // @[Breakpoint.scala 48:8:chipyard.TestHarness.RocketConfig.fir@249522.4]
  wire  _T_102; // @[Breakpoint.scala 85:32:chipyard.TestHarness.RocketConfig.fir@249523.4]
  wire  _T_106; // @[Breakpoint.scala 95:51:chipyard.TestHarness.RocketConfig.fir@249533.6]
  assign _T = ~io_status_debug; // @[Breakpoint.scala 31:35:chipyard.TestHarness.RocketConfig.fir@249421.4]
  assign _T_3 = {io_bp_0_control_m,1'h0,io_bp_0_control_s,io_bp_0_control_u}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@249424.4]
  assign _T_4 = _T_3 >> io_status_prv; // @[Breakpoint.scala 31:68:chipyard.TestHarness.RocketConfig.fir@249425.4]
  assign _T_6 = _T & _T_4[0]; // @[Breakpoint.scala 31:50:chipyard.TestHarness.RocketConfig.fir@249427.4]
  assign _T_7 = _T_6 & io_bp_0_control_r; // @[Breakpoint.scala 83:16:chipyard.TestHarness.RocketConfig.fir@249428.4]
  assign _T_9 = io_ea >= io_bp_0_address; // @[Breakpoint.scala 45:8:chipyard.TestHarness.RocketConfig.fir@249430.4]
  assign _T_11 = _T_9 ^ io_bp_0_control_tmatch[0]; // @[Breakpoint.scala 45:20:chipyard.TestHarness.RocketConfig.fir@249432.4]
  assign _T_12 = ~io_ea; // @[Breakpoint.scala 42:6:chipyard.TestHarness.RocketConfig.fir@249433.4]
  assign _T_15 = io_bp_0_control_tmatch[0] & io_bp_0_address[0]; // @[Breakpoint.scala 39:73:chipyard.TestHarness.RocketConfig.fir@249436.4]
  assign _T_17 = _T_15 & io_bp_0_address[1]; // @[Breakpoint.scala 39:73:chipyard.TestHarness.RocketConfig.fir@249438.4]
  assign _T_19 = _T_17 & io_bp_0_address[2]; // @[Breakpoint.scala 39:73:chipyard.TestHarness.RocketConfig.fir@249440.4]
  assign _T_22 = {_T_19,_T_17,_T_15,io_bp_0_control_tmatch[0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@249443.4]
  assign _GEN_11 = {{35'd0}, _T_22}; // @[Breakpoint.scala 42:9:chipyard.TestHarness.RocketConfig.fir@249444.4]
  assign _T_23 = _T_12 | _GEN_11; // @[Breakpoint.scala 42:9:chipyard.TestHarness.RocketConfig.fir@249444.4]
  assign _T_24 = ~io_bp_0_address; // @[Breakpoint.scala 42:24:chipyard.TestHarness.RocketConfig.fir@249445.4]
  assign _T_35 = _T_24 | _GEN_11; // @[Breakpoint.scala 42:33:chipyard.TestHarness.RocketConfig.fir@249456.4]
  assign _T_36 = _T_23 == _T_35; // @[Breakpoint.scala 42:19:chipyard.TestHarness.RocketConfig.fir@249457.4]
  assign _T_37 = io_bp_0_control_tmatch[1] ? _T_11 : _T_36; // @[Breakpoint.scala 48:8:chipyard.TestHarness.RocketConfig.fir@249458.4]
  assign _T_38 = _T_7 & _T_37; // @[Breakpoint.scala 83:32:chipyard.TestHarness.RocketConfig.fir@249459.4]
  assign _T_39 = _T_6 & io_bp_0_control_w; // @[Breakpoint.scala 84:16:chipyard.TestHarness.RocketConfig.fir@249460.4]
  assign _T_70 = _T_39 & _T_37; // @[Breakpoint.scala 84:32:chipyard.TestHarness.RocketConfig.fir@249491.4]
  assign _T_71 = _T_6 & io_bp_0_control_x; // @[Breakpoint.scala 85:16:chipyard.TestHarness.RocketConfig.fir@249492.4]
  assign _T_73 = io_pc >= io_bp_0_address; // @[Breakpoint.scala 45:8:chipyard.TestHarness.RocketConfig.fir@249494.4]
  assign _T_75 = _T_73 ^ io_bp_0_control_tmatch[0]; // @[Breakpoint.scala 45:20:chipyard.TestHarness.RocketConfig.fir@249496.4]
  assign _T_76 = ~io_pc; // @[Breakpoint.scala 42:6:chipyard.TestHarness.RocketConfig.fir@249497.4]
  assign _T_87 = _T_76 | _GEN_11; // @[Breakpoint.scala 42:9:chipyard.TestHarness.RocketConfig.fir@249508.4]
  assign _T_100 = _T_87 == _T_35; // @[Breakpoint.scala 42:19:chipyard.TestHarness.RocketConfig.fir@249521.4]
  assign _T_101 = io_bp_0_control_tmatch[1] ? _T_75 : _T_100; // @[Breakpoint.scala 48:8:chipyard.TestHarness.RocketConfig.fir@249522.4]
  assign _T_102 = _T_71 & _T_101; // @[Breakpoint.scala 85:32:chipyard.TestHarness.RocketConfig.fir@249523.4]
  assign _T_106 = ~io_bp_0_control_action; // @[Breakpoint.scala 95:51:chipyard.TestHarness.RocketConfig.fir@249533.6]
  assign io_xcpt_if = _T_102 & _T_106; // @[Breakpoint.scala 74:14:chipyard.TestHarness.RocketConfig.fir@249415.4 Breakpoint.scala 97:40:chipyard.TestHarness.RocketConfig.fir@249554.6]
  assign io_xcpt_ld = _T_38 & _T_106; // @[Breakpoint.scala 75:14:chipyard.TestHarness.RocketConfig.fir@249416.4 Breakpoint.scala 95:40:chipyard.TestHarness.RocketConfig.fir@249534.6]
  assign io_xcpt_st = _T_70 & _T_106; // @[Breakpoint.scala 76:14:chipyard.TestHarness.RocketConfig.fir@249417.4 Breakpoint.scala 96:40:chipyard.TestHarness.RocketConfig.fir@249544.6]
  assign io_debug_if = _T_102 & io_bp_0_control_action; // @[Breakpoint.scala 77:15:chipyard.TestHarness.RocketConfig.fir@249418.4 Breakpoint.scala 97:73:chipyard.TestHarness.RocketConfig.fir@249556.6]
  assign io_debug_ld = _T_38 & io_bp_0_control_action; // @[Breakpoint.scala 78:15:chipyard.TestHarness.RocketConfig.fir@249419.4 Breakpoint.scala 95:73:chipyard.TestHarness.RocketConfig.fir@249536.6]
  assign io_debug_st = _T_70 & io_bp_0_control_action; // @[Breakpoint.scala 79:15:chipyard.TestHarness.RocketConfig.fir@249420.4 Breakpoint.scala 96:73:chipyard.TestHarness.RocketConfig.fir@249546.6]
endmodule
