module RoundAnyRawFNToRecFN_3( // @[:chipyard.TestHarness.RocketConfig.fir@236253.2]
  input         io_invalidExc, // @[:chipyard.TestHarness.RocketConfig.fir@236254.4]
  input         io_in_isNaN, // @[:chipyard.TestHarness.RocketConfig.fir@236254.4]
  input         io_in_isInf, // @[:chipyard.TestHarness.RocketConfig.fir@236254.4]
  input         io_in_isZero, // @[:chipyard.TestHarness.RocketConfig.fir@236254.4]
  input         io_in_sign, // @[:chipyard.TestHarness.RocketConfig.fir@236254.4]
  input  [12:0] io_in_sExp, // @[:chipyard.TestHarness.RocketConfig.fir@236254.4]
  input  [53:0] io_in_sig, // @[:chipyard.TestHarness.RocketConfig.fir@236254.4]
  input  [2:0]  io_roundingMode, // @[:chipyard.TestHarness.RocketConfig.fir@236254.4]
  output [32:0] io_out, // @[:chipyard.TestHarness.RocketConfig.fir@236254.4]
  output [4:0]  io_exceptionFlags // @[:chipyard.TestHarness.RocketConfig.fir@236254.4]
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53:chipyard.TestHarness.RocketConfig.fir@236257.4]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53:chipyard.TestHarness.RocketConfig.fir@236259.4]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53:chipyard.TestHarness.RocketConfig.fir@236260.4]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53:chipyard.TestHarness.RocketConfig.fir@236261.4]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53:chipyard.TestHarness.RocketConfig.fir@236262.4]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27:chipyard.TestHarness.RocketConfig.fir@236263.4]
  wire  _T_1; // @[RoundAnyRawFNToRecFN.scala 96:66:chipyard.TestHarness.RocketConfig.fir@236264.4]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63:chipyard.TestHarness.RocketConfig.fir@236265.4]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42:chipyard.TestHarness.RocketConfig.fir@236266.4]
  wire [13:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 108:24:chipyard.TestHarness.RocketConfig.fir@236267.4]
  wire  _T_5; // @[RoundAnyRawFNToRecFN.scala 115:60:chipyard.TestHarness.RocketConfig.fir@236270.4]
  wire [26:0] adjustedSig; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236271.4]
  wire [8:0] _T_7; // @[primitives.scala 51:21:chipyard.TestHarness.RocketConfig.fir@236285.4]
  wire [64:0] _T_14; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@236292.4]
  wire [15:0] _T_20; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236298.4]
  wire [15:0] _T_22; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@236300.4]
  wire [15:0] _T_24; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@236302.4]
  wire [15:0] _T_25; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@236303.4]
  wire [15:0] _GEN_0; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236308.4]
  wire [15:0] _T_30; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236308.4]
  wire [15:0] _T_32; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@236310.4]
  wire [15:0] _T_34; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@236312.4]
  wire [15:0] _T_35; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@236313.4]
  wire [15:0] _GEN_1; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236318.4]
  wire [15:0] _T_40; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236318.4]
  wire [15:0] _T_42; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@236320.4]
  wire [15:0] _T_44; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@236322.4]
  wire [15:0] _T_45; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@236323.4]
  wire [15:0] _GEN_2; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236328.4]
  wire [15:0] _T_50; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236328.4]
  wire [15:0] _T_52; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@236330.4]
  wire [15:0] _T_54; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@236332.4]
  wire [15:0] _T_55; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@236333.4]
  wire [21:0] _T_72; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236350.4]
  wire [21:0] _T_73; // @[primitives.scala 74:36:chipyard.TestHarness.RocketConfig.fir@236351.4]
  wire [21:0] _T_74; // @[primitives.scala 74:21:chipyard.TestHarness.RocketConfig.fir@236352.4]
  wire [21:0] _T_75; // @[primitives.scala 74:17:chipyard.TestHarness.RocketConfig.fir@236353.4]
  wire [24:0] _T_76; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236354.4]
  wire [2:0] _T_86; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236364.4]
  wire [2:0] _T_87; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@236365.4]
  wire [24:0] _T_88; // @[primitives.scala 66:24:chipyard.TestHarness.RocketConfig.fir@236366.4]
  wire [24:0] _T_89; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@236367.4]
  wire [26:0] _T_91; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236369.4]
  wire [26:0] _T_93; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236371.4]
  wire [26:0] _T_94; // @[RoundAnyRawFNToRecFN.scala 161:28:chipyard.TestHarness.RocketConfig.fir@236372.4]
  wire [26:0] _T_95; // @[RoundAnyRawFNToRecFN.scala 161:46:chipyard.TestHarness.RocketConfig.fir@236373.4]
  wire [26:0] _T_96; // @[RoundAnyRawFNToRecFN.scala 162:40:chipyard.TestHarness.RocketConfig.fir@236374.4]
  wire  _T_97; // @[RoundAnyRawFNToRecFN.scala 162:56:chipyard.TestHarness.RocketConfig.fir@236375.4]
  wire [26:0] _T_98; // @[RoundAnyRawFNToRecFN.scala 163:42:chipyard.TestHarness.RocketConfig.fir@236376.4]
  wire  _T_99; // @[RoundAnyRawFNToRecFN.scala 163:62:chipyard.TestHarness.RocketConfig.fir@236377.4]
  wire  _T_100; // @[RoundAnyRawFNToRecFN.scala 164:36:chipyard.TestHarness.RocketConfig.fir@236378.4]
  wire  _T_101; // @[RoundAnyRawFNToRecFN.scala 167:38:chipyard.TestHarness.RocketConfig.fir@236379.4]
  wire  _T_102; // @[RoundAnyRawFNToRecFN.scala 167:67:chipyard.TestHarness.RocketConfig.fir@236380.4]
  wire  _T_103; // @[RoundAnyRawFNToRecFN.scala 169:29:chipyard.TestHarness.RocketConfig.fir@236381.4]
  wire  _T_104; // @[RoundAnyRawFNToRecFN.scala 168:31:chipyard.TestHarness.RocketConfig.fir@236382.4]
  wire [26:0] _T_105; // @[RoundAnyRawFNToRecFN.scala 172:32:chipyard.TestHarness.RocketConfig.fir@236383.4]
  wire [25:0] _T_107; // @[RoundAnyRawFNToRecFN.scala 172:49:chipyard.TestHarness.RocketConfig.fir@236385.4]
  wire  _T_108; // @[RoundAnyRawFNToRecFN.scala 173:49:chipyard.TestHarness.RocketConfig.fir@236386.4]
  wire  _T_109; // @[RoundAnyRawFNToRecFN.scala 174:30:chipyard.TestHarness.RocketConfig.fir@236387.4]
  wire  _T_110; // @[RoundAnyRawFNToRecFN.scala 173:64:chipyard.TestHarness.RocketConfig.fir@236388.4]
  wire [25:0] _T_112; // @[RoundAnyRawFNToRecFN.scala 173:25:chipyard.TestHarness.RocketConfig.fir@236390.4]
  wire [25:0] _T_113; // @[RoundAnyRawFNToRecFN.scala 173:21:chipyard.TestHarness.RocketConfig.fir@236391.4]
  wire [25:0] _T_114; // @[RoundAnyRawFNToRecFN.scala 172:61:chipyard.TestHarness.RocketConfig.fir@236392.4]
  wire [26:0] _T_115; // @[RoundAnyRawFNToRecFN.scala 178:32:chipyard.TestHarness.RocketConfig.fir@236393.4]
  wire [26:0] _T_116; // @[RoundAnyRawFNToRecFN.scala 178:30:chipyard.TestHarness.RocketConfig.fir@236394.4]
  wire  _T_118; // @[RoundAnyRawFNToRecFN.scala 179:42:chipyard.TestHarness.RocketConfig.fir@236396.4]
  wire [25:0] _T_120; // @[RoundAnyRawFNToRecFN.scala 179:24:chipyard.TestHarness.RocketConfig.fir@236398.4]
  wire [25:0] _GEN_3; // @[RoundAnyRawFNToRecFN.scala 178:47:chipyard.TestHarness.RocketConfig.fir@236399.4]
  wire [25:0] _T_121; // @[RoundAnyRawFNToRecFN.scala 178:47:chipyard.TestHarness.RocketConfig.fir@236399.4]
  wire [25:0] _T_122; // @[RoundAnyRawFNToRecFN.scala 171:16:chipyard.TestHarness.RocketConfig.fir@236400.4]
  wire [2:0] _T_124; // @[RoundAnyRawFNToRecFN.scala 183:69:chipyard.TestHarness.RocketConfig.fir@236402.4]
  wire [13:0] _GEN_4; // @[RoundAnyRawFNToRecFN.scala 183:40:chipyard.TestHarness.RocketConfig.fir@236403.4]
  wire [14:0] _T_125; // @[RoundAnyRawFNToRecFN.scala 183:40:chipyard.TestHarness.RocketConfig.fir@236403.4]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37:chipyard.TestHarness.RocketConfig.fir@236404.4]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 189:27:chipyard.TestHarness.RocketConfig.fir@236407.4]
  wire [7:0] _T_130; // @[RoundAnyRawFNToRecFN.scala 194:30:chipyard.TestHarness.RocketConfig.fir@236410.4]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50:chipyard.TestHarness.RocketConfig.fir@236411.4]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31:chipyard.TestHarness.RocketConfig.fir@236413.4]
  wire  _T_139; // @[RoundAnyRawFNToRecFN.scala 203:70:chipyard.TestHarness.RocketConfig.fir@236421.4]
  wire  _T_142; // @[RoundAnyRawFNToRecFN.scala 205:67:chipyard.TestHarness.RocketConfig.fir@236424.4]
  wire  _T_143; // @[RoundAnyRawFNToRecFN.scala 207:29:chipyard.TestHarness.RocketConfig.fir@236425.4]
  wire  _T_144; // @[RoundAnyRawFNToRecFN.scala 206:46:chipyard.TestHarness.RocketConfig.fir@236426.4]
  wire [5:0] _T_148; // @[RoundAnyRawFNToRecFN.scala 218:48:chipyard.TestHarness.RocketConfig.fir@236430.4]
  wire  _T_149; // @[RoundAnyRawFNToRecFN.scala 218:62:chipyard.TestHarness.RocketConfig.fir@236431.4]
  wire  _T_150; // @[RoundAnyRawFNToRecFN.scala 218:32:chipyard.TestHarness.RocketConfig.fir@236432.4]
  wire  _T_154; // @[RoundAnyRawFNToRecFN.scala 218:74:chipyard.TestHarness.RocketConfig.fir@236436.4]
  wire  _T_159; // @[RoundAnyRawFNToRecFN.scala 221:34:chipyard.TestHarness.RocketConfig.fir@236441.4]
  wire  _T_161; // @[RoundAnyRawFNToRecFN.scala 224:38:chipyard.TestHarness.RocketConfig.fir@236443.4]
  wire  _T_162; // @[RoundAnyRawFNToRecFN.scala 225:45:chipyard.TestHarness.RocketConfig.fir@236444.4]
  wire  _T_163; // @[RoundAnyRawFNToRecFN.scala 225:60:chipyard.TestHarness.RocketConfig.fir@236445.4]
  wire  _T_164; // @[RoundAnyRawFNToRecFN.scala 220:27:chipyard.TestHarness.RocketConfig.fir@236446.4]
  wire  _T_165; // @[RoundAnyRawFNToRecFN.scala 219:76:chipyard.TestHarness.RocketConfig.fir@236447.4]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40:chipyard.TestHarness.RocketConfig.fir@236448.4]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49:chipyard.TestHarness.RocketConfig.fir@236450.4]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34:chipyard.TestHarness.RocketConfig.fir@236452.4]
  wire  _T_168; // @[RoundAnyRawFNToRecFN.scala 235:22:chipyard.TestHarness.RocketConfig.fir@236454.4]
  wire  _T_169; // @[RoundAnyRawFNToRecFN.scala 235:36:chipyard.TestHarness.RocketConfig.fir@236455.4]
  wire  _T_170; // @[RoundAnyRawFNToRecFN.scala 235:33:chipyard.TestHarness.RocketConfig.fir@236456.4]
  wire  _T_171; // @[RoundAnyRawFNToRecFN.scala 235:64:chipyard.TestHarness.RocketConfig.fir@236457.4]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61:chipyard.TestHarness.RocketConfig.fir@236458.4]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32:chipyard.TestHarness.RocketConfig.fir@236459.4]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32:chipyard.TestHarness.RocketConfig.fir@236460.4]
  wire  _T_172; // @[RoundAnyRawFNToRecFN.scala 238:43:chipyard.TestHarness.RocketConfig.fir@236461.4]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28:chipyard.TestHarness.RocketConfig.fir@236462.4]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60:chipyard.TestHarness.RocketConfig.fir@236464.4]
  wire  _T_174; // @[RoundAnyRawFNToRecFN.scala 243:20:chipyard.TestHarness.RocketConfig.fir@236465.4]
  wire  _T_175; // @[RoundAnyRawFNToRecFN.scala 243:60:chipyard.TestHarness.RocketConfig.fir@236466.4]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45:chipyard.TestHarness.RocketConfig.fir@236467.4]
  wire  _T_176; // @[RoundAnyRawFNToRecFN.scala 244:42:chipyard.TestHarness.RocketConfig.fir@236468.4]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39:chipyard.TestHarness.RocketConfig.fir@236469.4]
  wire  _T_177; // @[RoundAnyRawFNToRecFN.scala 246:45:chipyard.TestHarness.RocketConfig.fir@236470.4]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32:chipyard.TestHarness.RocketConfig.fir@236471.4]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22:chipyard.TestHarness.RocketConfig.fir@236472.4]
  wire  _T_178; // @[RoundAnyRawFNToRecFN.scala 251:32:chipyard.TestHarness.RocketConfig.fir@236473.4]
  wire [8:0] _T_179; // @[RoundAnyRawFNToRecFN.scala 251:18:chipyard.TestHarness.RocketConfig.fir@236474.4]
  wire [8:0] _T_180; // @[RoundAnyRawFNToRecFN.scala 251:14:chipyard.TestHarness.RocketConfig.fir@236475.4]
  wire [8:0] _T_181; // @[RoundAnyRawFNToRecFN.scala 250:24:chipyard.TestHarness.RocketConfig.fir@236476.4]
  wire [8:0] _T_183; // @[RoundAnyRawFNToRecFN.scala 255:18:chipyard.TestHarness.RocketConfig.fir@236478.4]
  wire [8:0] _T_184; // @[RoundAnyRawFNToRecFN.scala 255:14:chipyard.TestHarness.RocketConfig.fir@236479.4]
  wire [8:0] _T_185; // @[RoundAnyRawFNToRecFN.scala 254:17:chipyard.TestHarness.RocketConfig.fir@236480.4]
  wire [8:0] _T_186; // @[RoundAnyRawFNToRecFN.scala 259:18:chipyard.TestHarness.RocketConfig.fir@236481.4]
  wire [8:0] _T_187; // @[RoundAnyRawFNToRecFN.scala 259:14:chipyard.TestHarness.RocketConfig.fir@236482.4]
  wire [8:0] _T_188; // @[RoundAnyRawFNToRecFN.scala 258:17:chipyard.TestHarness.RocketConfig.fir@236483.4]
  wire [8:0] _T_189; // @[RoundAnyRawFNToRecFN.scala 263:18:chipyard.TestHarness.RocketConfig.fir@236484.4]
  wire [8:0] _T_190; // @[RoundAnyRawFNToRecFN.scala 263:14:chipyard.TestHarness.RocketConfig.fir@236485.4]
  wire [8:0] _T_191; // @[RoundAnyRawFNToRecFN.scala 262:17:chipyard.TestHarness.RocketConfig.fir@236486.4]
  wire [8:0] _T_192; // @[RoundAnyRawFNToRecFN.scala 267:16:chipyard.TestHarness.RocketConfig.fir@236487.4]
  wire [8:0] _T_193; // @[RoundAnyRawFNToRecFN.scala 266:18:chipyard.TestHarness.RocketConfig.fir@236488.4]
  wire [8:0] _T_194; // @[RoundAnyRawFNToRecFN.scala 271:16:chipyard.TestHarness.RocketConfig.fir@236489.4]
  wire [8:0] _T_195; // @[RoundAnyRawFNToRecFN.scala 270:15:chipyard.TestHarness.RocketConfig.fir@236490.4]
  wire [8:0] _T_196; // @[RoundAnyRawFNToRecFN.scala 275:16:chipyard.TestHarness.RocketConfig.fir@236491.4]
  wire [8:0] _T_197; // @[RoundAnyRawFNToRecFN.scala 274:15:chipyard.TestHarness.RocketConfig.fir@236492.4]
  wire [8:0] _T_198; // @[RoundAnyRawFNToRecFN.scala 276:16:chipyard.TestHarness.RocketConfig.fir@236493.4]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77:chipyard.TestHarness.RocketConfig.fir@236494.4]
  wire  _T_199; // @[RoundAnyRawFNToRecFN.scala 278:22:chipyard.TestHarness.RocketConfig.fir@236495.4]
  wire  _T_200; // @[RoundAnyRawFNToRecFN.scala 278:38:chipyard.TestHarness.RocketConfig.fir@236496.4]
  wire [22:0] _T_201; // @[RoundAnyRawFNToRecFN.scala 279:16:chipyard.TestHarness.RocketConfig.fir@236497.4]
  wire [22:0] _T_202; // @[RoundAnyRawFNToRecFN.scala 278:12:chipyard.TestHarness.RocketConfig.fir@236498.4]
  wire [22:0] _T_204; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@236500.4]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11:chipyard.TestHarness.RocketConfig.fir@236501.4]
  wire [9:0] _T_205; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236502.4]
  wire [1:0] _T_207; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236505.4]
  wire [2:0] _T_209; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236507.4]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53:chipyard.TestHarness.RocketConfig.fir@236257.4]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53:chipyard.TestHarness.RocketConfig.fir@236259.4]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53:chipyard.TestHarness.RocketConfig.fir@236260.4]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53:chipyard.TestHarness.RocketConfig.fir@236261.4]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53:chipyard.TestHarness.RocketConfig.fir@236262.4]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27:chipyard.TestHarness.RocketConfig.fir@236263.4]
  assign _T_1 = ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:66:chipyard.TestHarness.RocketConfig.fir@236264.4]
  assign _T_2 = roundingMode_max & _T_1; // @[RoundAnyRawFNToRecFN.scala 96:63:chipyard.TestHarness.RocketConfig.fir@236265.4]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42:chipyard.TestHarness.RocketConfig.fir@236266.4]
  assign sAdjustedExp = $signed(io_in_sExp) - 13'sh700; // @[RoundAnyRawFNToRecFN.scala 108:24:chipyard.TestHarness.RocketConfig.fir@236267.4]
  assign _T_5 = |io_in_sig[27:0]; // @[RoundAnyRawFNToRecFN.scala 115:60:chipyard.TestHarness.RocketConfig.fir@236270.4]
  assign adjustedSig = {io_in_sig[53:28],_T_5}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236271.4]
  assign _T_7 = ~sAdjustedExp[8:0]; // @[primitives.scala 51:21:chipyard.TestHarness.RocketConfig.fir@236285.4]
  assign _T_14 = -65'sh10000000000000000 >>> _T_7[5:0]; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@236292.4]
  assign _T_20 = {{8'd0}, _T_14[57:50]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236298.4]
  assign _T_22 = {_T_14[49:42], 8'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@236300.4]
  assign _T_24 = _T_22 & 16'hff00; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@236302.4]
  assign _T_25 = _T_20 | _T_24; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@236303.4]
  assign _GEN_0 = {{4'd0}, _T_25[15:4]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236308.4]
  assign _T_30 = _GEN_0 & 16'hf0f; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236308.4]
  assign _T_32 = {_T_25[11:0], 4'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@236310.4]
  assign _T_34 = _T_32 & 16'hf0f0; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@236312.4]
  assign _T_35 = _T_30 | _T_34; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@236313.4]
  assign _GEN_1 = {{2'd0}, _T_35[15:2]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236318.4]
  assign _T_40 = _GEN_1 & 16'h3333; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236318.4]
  assign _T_42 = {_T_35[13:0], 2'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@236320.4]
  assign _T_44 = _T_42 & 16'hcccc; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@236322.4]
  assign _T_45 = _T_40 | _T_44; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@236323.4]
  assign _GEN_2 = {{1'd0}, _T_45[15:1]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236328.4]
  assign _T_50 = _GEN_2 & 16'h5555; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@236328.4]
  assign _T_52 = {_T_45[14:0], 1'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@236330.4]
  assign _T_54 = _T_52 & 16'haaaa; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@236332.4]
  assign _T_55 = _T_50 | _T_54; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@236333.4]
  assign _T_72 = {_T_55,_T_14[58],_T_14[59],_T_14[60],_T_14[61],_T_14[62],_T_14[63]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236350.4]
  assign _T_73 = ~_T_72; // @[primitives.scala 74:36:chipyard.TestHarness.RocketConfig.fir@236351.4]
  assign _T_74 = _T_7[6] ? 22'h0 : _T_73; // @[primitives.scala 74:21:chipyard.TestHarness.RocketConfig.fir@236352.4]
  assign _T_75 = ~_T_74; // @[primitives.scala 74:17:chipyard.TestHarness.RocketConfig.fir@236353.4]
  assign _T_76 = {_T_75,3'h7}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236354.4]
  assign _T_86 = {_T_14[0],_T_14[1],_T_14[2]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236364.4]
  assign _T_87 = _T_7[6] ? _T_86 : 3'h0; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@236365.4]
  assign _T_88 = _T_7[7] ? _T_76 : {{22'd0}, _T_87}; // @[primitives.scala 66:24:chipyard.TestHarness.RocketConfig.fir@236366.4]
  assign _T_89 = _T_7[8] ? _T_88 : 25'h0; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@236367.4]
  assign _T_91 = {_T_89,2'h3}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236369.4]
  assign _T_93 = {1'h0,_T_91[26:1]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236371.4]
  assign _T_94 = ~_T_93; // @[RoundAnyRawFNToRecFN.scala 161:28:chipyard.TestHarness.RocketConfig.fir@236372.4]
  assign _T_95 = _T_94 & _T_91; // @[RoundAnyRawFNToRecFN.scala 161:46:chipyard.TestHarness.RocketConfig.fir@236373.4]
  assign _T_96 = adjustedSig & _T_95; // @[RoundAnyRawFNToRecFN.scala 162:40:chipyard.TestHarness.RocketConfig.fir@236374.4]
  assign _T_97 = |_T_96; // @[RoundAnyRawFNToRecFN.scala 162:56:chipyard.TestHarness.RocketConfig.fir@236375.4]
  assign _T_98 = adjustedSig & _T_93; // @[RoundAnyRawFNToRecFN.scala 163:42:chipyard.TestHarness.RocketConfig.fir@236376.4]
  assign _T_99 = |_T_98; // @[RoundAnyRawFNToRecFN.scala 163:62:chipyard.TestHarness.RocketConfig.fir@236377.4]
  assign _T_100 = _T_97 | _T_99; // @[RoundAnyRawFNToRecFN.scala 164:36:chipyard.TestHarness.RocketConfig.fir@236378.4]
  assign _T_101 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38:chipyard.TestHarness.RocketConfig.fir@236379.4]
  assign _T_102 = _T_101 & _T_97; // @[RoundAnyRawFNToRecFN.scala 167:67:chipyard.TestHarness.RocketConfig.fir@236380.4]
  assign _T_103 = roundMagUp & _T_100; // @[RoundAnyRawFNToRecFN.scala 169:29:chipyard.TestHarness.RocketConfig.fir@236381.4]
  assign _T_104 = _T_102 | _T_103; // @[RoundAnyRawFNToRecFN.scala 168:31:chipyard.TestHarness.RocketConfig.fir@236382.4]
  assign _T_105 = adjustedSig | _T_91; // @[RoundAnyRawFNToRecFN.scala 172:32:chipyard.TestHarness.RocketConfig.fir@236383.4]
  assign _T_107 = _T_105[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49:chipyard.TestHarness.RocketConfig.fir@236385.4]
  assign _T_108 = roundingMode_near_even & _T_97; // @[RoundAnyRawFNToRecFN.scala 173:49:chipyard.TestHarness.RocketConfig.fir@236386.4]
  assign _T_109 = ~_T_99; // @[RoundAnyRawFNToRecFN.scala 174:30:chipyard.TestHarness.RocketConfig.fir@236387.4]
  assign _T_110 = _T_108 & _T_109; // @[RoundAnyRawFNToRecFN.scala 173:64:chipyard.TestHarness.RocketConfig.fir@236388.4]
  assign _T_112 = _T_110 ? _T_91[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25:chipyard.TestHarness.RocketConfig.fir@236390.4]
  assign _T_113 = ~_T_112; // @[RoundAnyRawFNToRecFN.scala 173:21:chipyard.TestHarness.RocketConfig.fir@236391.4]
  assign _T_114 = _T_107 & _T_113; // @[RoundAnyRawFNToRecFN.scala 172:61:chipyard.TestHarness.RocketConfig.fir@236392.4]
  assign _T_115 = ~_T_91; // @[RoundAnyRawFNToRecFN.scala 178:32:chipyard.TestHarness.RocketConfig.fir@236393.4]
  assign _T_116 = adjustedSig & _T_115; // @[RoundAnyRawFNToRecFN.scala 178:30:chipyard.TestHarness.RocketConfig.fir@236394.4]
  assign _T_118 = roundingMode_odd & _T_100; // @[RoundAnyRawFNToRecFN.scala 179:42:chipyard.TestHarness.RocketConfig.fir@236396.4]
  assign _T_120 = _T_118 ? _T_95[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 179:24:chipyard.TestHarness.RocketConfig.fir@236398.4]
  assign _GEN_3 = {{1'd0}, _T_116[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47:chipyard.TestHarness.RocketConfig.fir@236399.4]
  assign _T_121 = _GEN_3 | _T_120; // @[RoundAnyRawFNToRecFN.scala 178:47:chipyard.TestHarness.RocketConfig.fir@236399.4]
  assign _T_122 = _T_104 ? _T_114 : _T_121; // @[RoundAnyRawFNToRecFN.scala 171:16:chipyard.TestHarness.RocketConfig.fir@236400.4]
  assign _T_124 = {1'b0,$signed(_T_122[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69:chipyard.TestHarness.RocketConfig.fir@236402.4]
  assign _GEN_4 = {{11{_T_124[2]}},_T_124}; // @[RoundAnyRawFNToRecFN.scala 183:40:chipyard.TestHarness.RocketConfig.fir@236403.4]
  assign _T_125 = $signed(sAdjustedExp) + $signed(_GEN_4); // @[RoundAnyRawFNToRecFN.scala 183:40:chipyard.TestHarness.RocketConfig.fir@236403.4]
  assign common_expOut = _T_125[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37:chipyard.TestHarness.RocketConfig.fir@236404.4]
  assign common_fractOut = _T_122[22:0]; // @[RoundAnyRawFNToRecFN.scala 189:27:chipyard.TestHarness.RocketConfig.fir@236407.4]
  assign _T_130 = _T_125[14:7]; // @[RoundAnyRawFNToRecFN.scala 194:30:chipyard.TestHarness.RocketConfig.fir@236410.4]
  assign common_overflow = $signed(_T_130) >= 8'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50:chipyard.TestHarness.RocketConfig.fir@236411.4]
  assign common_totalUnderflow = $signed(_T_125) < 15'sh6b; // @[RoundAnyRawFNToRecFN.scala 198:31:chipyard.TestHarness.RocketConfig.fir@236413.4]
  assign _T_139 = |adjustedSig[1:0]; // @[RoundAnyRawFNToRecFN.scala 203:70:chipyard.TestHarness.RocketConfig.fir@236421.4]
  assign _T_142 = _T_101 & adjustedSig[1]; // @[RoundAnyRawFNToRecFN.scala 205:67:chipyard.TestHarness.RocketConfig.fir@236424.4]
  assign _T_143 = roundMagUp & _T_139; // @[RoundAnyRawFNToRecFN.scala 207:29:chipyard.TestHarness.RocketConfig.fir@236425.4]
  assign _T_144 = _T_142 | _T_143; // @[RoundAnyRawFNToRecFN.scala 206:46:chipyard.TestHarness.RocketConfig.fir@236426.4]
  assign _T_148 = sAdjustedExp[13:8]; // @[RoundAnyRawFNToRecFN.scala 218:48:chipyard.TestHarness.RocketConfig.fir@236430.4]
  assign _T_149 = $signed(_T_148) <= 6'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62:chipyard.TestHarness.RocketConfig.fir@236431.4]
  assign _T_150 = _T_100 & _T_149; // @[RoundAnyRawFNToRecFN.scala 218:32:chipyard.TestHarness.RocketConfig.fir@236432.4]
  assign _T_154 = _T_150 & _T_91[2]; // @[RoundAnyRawFNToRecFN.scala 218:74:chipyard.TestHarness.RocketConfig.fir@236436.4]
  assign _T_159 = ~_T_91[3]; // @[RoundAnyRawFNToRecFN.scala 221:34:chipyard.TestHarness.RocketConfig.fir@236441.4]
  assign _T_161 = _T_159 & _T_122[24]; // @[RoundAnyRawFNToRecFN.scala 224:38:chipyard.TestHarness.RocketConfig.fir@236443.4]
  assign _T_162 = _T_161 & _T_97; // @[RoundAnyRawFNToRecFN.scala 225:45:chipyard.TestHarness.RocketConfig.fir@236444.4]
  assign _T_163 = _T_162 & _T_144; // @[RoundAnyRawFNToRecFN.scala 225:60:chipyard.TestHarness.RocketConfig.fir@236445.4]
  assign _T_164 = ~_T_163; // @[RoundAnyRawFNToRecFN.scala 220:27:chipyard.TestHarness.RocketConfig.fir@236446.4]
  assign _T_165 = _T_154 & _T_164; // @[RoundAnyRawFNToRecFN.scala 219:76:chipyard.TestHarness.RocketConfig.fir@236447.4]
  assign common_underflow = common_totalUnderflow | _T_165; // @[RoundAnyRawFNToRecFN.scala 215:40:chipyard.TestHarness.RocketConfig.fir@236448.4]
  assign common_inexact = common_totalUnderflow | _T_100; // @[RoundAnyRawFNToRecFN.scala 228:49:chipyard.TestHarness.RocketConfig.fir@236450.4]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34:chipyard.TestHarness.RocketConfig.fir@236452.4]
  assign _T_168 = ~isNaNOut; // @[RoundAnyRawFNToRecFN.scala 235:22:chipyard.TestHarness.RocketConfig.fir@236454.4]
  assign _T_169 = ~io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 235:36:chipyard.TestHarness.RocketConfig.fir@236455.4]
  assign _T_170 = _T_168 & _T_169; // @[RoundAnyRawFNToRecFN.scala 235:33:chipyard.TestHarness.RocketConfig.fir@236456.4]
  assign _T_171 = ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:64:chipyard.TestHarness.RocketConfig.fir@236457.4]
  assign commonCase = _T_170 & _T_171; // @[RoundAnyRawFNToRecFN.scala 235:61:chipyard.TestHarness.RocketConfig.fir@236458.4]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32:chipyard.TestHarness.RocketConfig.fir@236459.4]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32:chipyard.TestHarness.RocketConfig.fir@236460.4]
  assign _T_172 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43:chipyard.TestHarness.RocketConfig.fir@236461.4]
  assign inexact = overflow | _T_172; // @[RoundAnyRawFNToRecFN.scala 238:28:chipyard.TestHarness.RocketConfig.fir@236462.4]
  assign overflow_roundMagUp = _T_101 | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60:chipyard.TestHarness.RocketConfig.fir@236464.4]
  assign _T_174 = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20:chipyard.TestHarness.RocketConfig.fir@236465.4]
  assign _T_175 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60:chipyard.TestHarness.RocketConfig.fir@236466.4]
  assign pegMinNonzeroMagOut = _T_174 & _T_175; // @[RoundAnyRawFNToRecFN.scala 243:45:chipyard.TestHarness.RocketConfig.fir@236467.4]
  assign _T_176 = ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:42:chipyard.TestHarness.RocketConfig.fir@236468.4]
  assign pegMaxFiniteMagOut = overflow & _T_176; // @[RoundAnyRawFNToRecFN.scala 244:39:chipyard.TestHarness.RocketConfig.fir@236469.4]
  assign _T_177 = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45:chipyard.TestHarness.RocketConfig.fir@236470.4]
  assign notNaN_isInfOut = io_in_isInf | _T_177; // @[RoundAnyRawFNToRecFN.scala 246:32:chipyard.TestHarness.RocketConfig.fir@236471.4]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22:chipyard.TestHarness.RocketConfig.fir@236472.4]
  assign _T_178 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32:chipyard.TestHarness.RocketConfig.fir@236473.4]
  assign _T_179 = _T_178 ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18:chipyard.TestHarness.RocketConfig.fir@236474.4]
  assign _T_180 = ~_T_179; // @[RoundAnyRawFNToRecFN.scala 251:14:chipyard.TestHarness.RocketConfig.fir@236475.4]
  assign _T_181 = common_expOut & _T_180; // @[RoundAnyRawFNToRecFN.scala 250:24:chipyard.TestHarness.RocketConfig.fir@236476.4]
  assign _T_183 = pegMinNonzeroMagOut ? 9'h194 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 255:18:chipyard.TestHarness.RocketConfig.fir@236478.4]
  assign _T_184 = ~_T_183; // @[RoundAnyRawFNToRecFN.scala 255:14:chipyard.TestHarness.RocketConfig.fir@236479.4]
  assign _T_185 = _T_181 & _T_184; // @[RoundAnyRawFNToRecFN.scala 254:17:chipyard.TestHarness.RocketConfig.fir@236480.4]
  assign _T_186 = pegMaxFiniteMagOut ? 9'h80 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 259:18:chipyard.TestHarness.RocketConfig.fir@236481.4]
  assign _T_187 = ~_T_186; // @[RoundAnyRawFNToRecFN.scala 259:14:chipyard.TestHarness.RocketConfig.fir@236482.4]
  assign _T_188 = _T_185 & _T_187; // @[RoundAnyRawFNToRecFN.scala 258:17:chipyard.TestHarness.RocketConfig.fir@236483.4]
  assign _T_189 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 263:18:chipyard.TestHarness.RocketConfig.fir@236484.4]
  assign _T_190 = ~_T_189; // @[RoundAnyRawFNToRecFN.scala 263:14:chipyard.TestHarness.RocketConfig.fir@236485.4]
  assign _T_191 = _T_188 & _T_190; // @[RoundAnyRawFNToRecFN.scala 262:17:chipyard.TestHarness.RocketConfig.fir@236486.4]
  assign _T_192 = pegMinNonzeroMagOut ? 9'h6b : 9'h0; // @[RoundAnyRawFNToRecFN.scala 267:16:chipyard.TestHarness.RocketConfig.fir@236487.4]
  assign _T_193 = _T_191 | _T_192; // @[RoundAnyRawFNToRecFN.scala 266:18:chipyard.TestHarness.RocketConfig.fir@236488.4]
  assign _T_194 = pegMaxFiniteMagOut ? 9'h17f : 9'h0; // @[RoundAnyRawFNToRecFN.scala 271:16:chipyard.TestHarness.RocketConfig.fir@236489.4]
  assign _T_195 = _T_193 | _T_194; // @[RoundAnyRawFNToRecFN.scala 270:15:chipyard.TestHarness.RocketConfig.fir@236490.4]
  assign _T_196 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 275:16:chipyard.TestHarness.RocketConfig.fir@236491.4]
  assign _T_197 = _T_195 | _T_196; // @[RoundAnyRawFNToRecFN.scala 274:15:chipyard.TestHarness.RocketConfig.fir@236492.4]
  assign _T_198 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 276:16:chipyard.TestHarness.RocketConfig.fir@236493.4]
  assign expOut = _T_197 | _T_198; // @[RoundAnyRawFNToRecFN.scala 275:77:chipyard.TestHarness.RocketConfig.fir@236494.4]
  assign _T_199 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22:chipyard.TestHarness.RocketConfig.fir@236495.4]
  assign _T_200 = _T_199 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38:chipyard.TestHarness.RocketConfig.fir@236496.4]
  assign _T_201 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 279:16:chipyard.TestHarness.RocketConfig.fir@236497.4]
  assign _T_202 = _T_200 ? _T_201 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12:chipyard.TestHarness.RocketConfig.fir@236498.4]
  assign _T_204 = pegMaxFiniteMagOut ? 23'h7fffff : 23'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@236500.4]
  assign fractOut = _T_202 | _T_204; // @[RoundAnyRawFNToRecFN.scala 281:11:chipyard.TestHarness.RocketConfig.fir@236501.4]
  assign _T_205 = {signOut,expOut}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236502.4]
  assign _T_207 = {underflow,inexact}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236505.4]
  assign _T_209 = {io_invalidExc,1'h0,overflow}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@236507.4]
  assign io_out = {_T_205,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12:chipyard.TestHarness.RocketConfig.fir@236504.4]
  assign io_exceptionFlags = {_T_209,_T_207}; // @[RoundAnyRawFNToRecFN.scala 285:23:chipyard.TestHarness.RocketConfig.fir@236509.4]
endmodule
