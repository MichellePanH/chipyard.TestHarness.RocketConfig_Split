module ClockGroupAggregator_1( // @[:chipyard.TestHarness.RocketConfig.fir@20914.2]
  input   auto_in_member_0_clock, // @[:chipyard.TestHarness.RocketConfig.fir@20915.4]
  input   auto_in_member_0_reset, // @[:chipyard.TestHarness.RocketConfig.fir@20915.4]
  output  auto_out_member_0_clock, // @[:chipyard.TestHarness.RocketConfig.fir@20915.4]
  output  auto_out_member_0_reset // @[:chipyard.TestHarness.RocketConfig.fir@20915.4]
);
  assign auto_out_member_0_clock = auto_in_member_0_clock; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@20929.4]
  assign auto_out_member_0_reset = auto_in_member_0_reset; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@20929.4]
endmodule
