module SimpleClockGroupSource( // @[:chipyard.TestHarness.RocketConfig.fir@19.2]
  input   clock, // @[:chipyard.TestHarness.RocketConfig.fir@20.4]
  input   reset, // @[:chipyard.TestHarness.RocketConfig.fir@21.4]
  output  auto_out_member_5_clock, // @[:chipyard.TestHarness.RocketConfig.fir@22.4]
  output  auto_out_member_5_reset, // @[:chipyard.TestHarness.RocketConfig.fir@22.4]
  output  auto_out_member_4_clock, // @[:chipyard.TestHarness.RocketConfig.fir@22.4]
  output  auto_out_member_4_reset, // @[:chipyard.TestHarness.RocketConfig.fir@22.4]
  output  auto_out_member_3_clock, // @[:chipyard.TestHarness.RocketConfig.fir@22.4]
  output  auto_out_member_3_reset, // @[:chipyard.TestHarness.RocketConfig.fir@22.4]
  output  auto_out_member_2_clock, // @[:chipyard.TestHarness.RocketConfig.fir@22.4]
  output  auto_out_member_2_reset, // @[:chipyard.TestHarness.RocketConfig.fir@22.4]
  output  auto_out_member_1_clock, // @[:chipyard.TestHarness.RocketConfig.fir@22.4]
  output  auto_out_member_1_reset, // @[:chipyard.TestHarness.RocketConfig.fir@22.4]
  output  auto_out_member_0_clock, // @[:chipyard.TestHarness.RocketConfig.fir@22.4]
  output  auto_out_member_0_reset // @[:chipyard.TestHarness.RocketConfig.fir@22.4]
);
  assign auto_out_member_5_clock = clock; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@29.4]
  assign auto_out_member_5_reset = reset; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@29.4]
  assign auto_out_member_4_clock = clock; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@29.4]
  assign auto_out_member_4_reset = reset; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@29.4]
  assign auto_out_member_3_clock = clock; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@29.4]
  assign auto_out_member_3_reset = reset; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@29.4]
  assign auto_out_member_2_clock = clock; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@29.4]
  assign auto_out_member_2_reset = reset; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@29.4]
  assign auto_out_member_1_clock = clock; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@29.4]
  assign auto_out_member_1_reset = reset; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@29.4]
  assign auto_out_member_0_clock = clock; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@29.4]
  assign auto_out_member_0_reset = reset; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@29.4]
endmodule
