module Arbiter( // @[:chipyard.TestHarness.RocketConfig.fir@240824.2]
  output        io_in_0_ready, // @[:chipyard.TestHarness.RocketConfig.fir@240827.4]
  input         io_in_0_valid, // @[:chipyard.TestHarness.RocketConfig.fir@240827.4]
  input  [26:0] io_in_0_bits_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@240827.4]
  output        io_in_1_ready, // @[:chipyard.TestHarness.RocketConfig.fir@240827.4]
  input         io_in_1_valid, // @[:chipyard.TestHarness.RocketConfig.fir@240827.4]
  input         io_in_1_bits_valid, // @[:chipyard.TestHarness.RocketConfig.fir@240827.4]
  input  [26:0] io_in_1_bits_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@240827.4]
  input         io_out_ready, // @[:chipyard.TestHarness.RocketConfig.fir@240827.4]
  output        io_out_valid, // @[:chipyard.TestHarness.RocketConfig.fir@240827.4]
  output        io_out_bits_valid, // @[:chipyard.TestHarness.RocketConfig.fir@240827.4]
  output [26:0] io_out_bits_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@240827.4]
  output        io_chosen // @[:chipyard.TestHarness.RocketConfig.fir@240827.4]
);
  wire  grant_1; // @[Arbiter.scala 31:78:chipyard.TestHarness.RocketConfig.fir@240837.4]
  wire  _T_2; // @[Arbiter.scala 135:19:chipyard.TestHarness.RocketConfig.fir@240842.4]
  assign grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78:chipyard.TestHarness.RocketConfig.fir@240837.4]
  assign _T_2 = ~grant_1; // @[Arbiter.scala 135:19:chipyard.TestHarness.RocketConfig.fir@240842.4]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14:chipyard.TestHarness.RocketConfig.fir@240839.4]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14:chipyard.TestHarness.RocketConfig.fir@240841.4]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16:chipyard.TestHarness.RocketConfig.fir@240844.4]
  assign io_out_bits_valid = io_in_0_valid | io_in_1_bits_valid; // @[Arbiter.scala 124:15:chipyard.TestHarness.RocketConfig.fir@240831.4 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@240835.6]
  assign io_out_bits_bits_addr = io_in_0_valid ? io_in_0_bits_bits_addr : io_in_1_bits_bits_addr; // @[Arbiter.scala 124:15:chipyard.TestHarness.RocketConfig.fir@240830.4 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@240834.6]
  assign io_chosen = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 123:13:chipyard.TestHarness.RocketConfig.fir@240829.4 Arbiter.scala 127:17:chipyard.TestHarness.RocketConfig.fir@240833.6]
endmodule
