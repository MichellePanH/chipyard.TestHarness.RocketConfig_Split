module DMIToTL( // @[:chipyard.TestHarness.RocketConfig.fir@126677.2]
  input         auto_out_a_ready, // @[:chipyard.TestHarness.RocketConfig.fir@126680.4]
  output        auto_out_a_valid, // @[:chipyard.TestHarness.RocketConfig.fir@126680.4]
  output [2:0]  auto_out_a_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@126680.4]
  output [8:0]  auto_out_a_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@126680.4]
  output [3:0]  auto_out_a_bits_mask, // @[:chipyard.TestHarness.RocketConfig.fir@126680.4]
  output [31:0] auto_out_a_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@126680.4]
  output        auto_out_d_ready, // @[:chipyard.TestHarness.RocketConfig.fir@126680.4]
  input         auto_out_d_valid, // @[:chipyard.TestHarness.RocketConfig.fir@126680.4]
  input         auto_out_d_bits_denied, // @[:chipyard.TestHarness.RocketConfig.fir@126680.4]
  input  [31:0] auto_out_d_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@126680.4]
  input         auto_out_d_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@126680.4]
  output        io_dmi_req_ready, // @[:chipyard.TestHarness.RocketConfig.fir@126681.4]
  input         io_dmi_req_valid, // @[:chipyard.TestHarness.RocketConfig.fir@126681.4]
  input  [6:0]  io_dmi_req_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@126681.4]
  input  [31:0] io_dmi_req_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@126681.4]
  input  [1:0]  io_dmi_req_bits_op, // @[:chipyard.TestHarness.RocketConfig.fir@126681.4]
  input         io_dmi_resp_ready, // @[:chipyard.TestHarness.RocketConfig.fir@126681.4]
  output        io_dmi_resp_valid, // @[:chipyard.TestHarness.RocketConfig.fir@126681.4]
  output [31:0] io_dmi_resp_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@126681.4]
  output [1:0]  io_dmi_resp_bits_resp // @[:chipyard.TestHarness.RocketConfig.fir@126681.4]
);
  wire [8:0] addr; // @[DMI.scala 97:46:chipyard.TestHarness.RocketConfig.fir@126692.4]
  wire  _T_100; // @[DMI.scala 111:30:chipyard.TestHarness.RocketConfig.fir@126824.4]
  wire  _T_101; // @[DMI.scala 112:37:chipyard.TestHarness.RocketConfig.fir@126836.6]
  wire [3:0] _GEN_2; // @[DMI.scala 112:64:chipyard.TestHarness.RocketConfig.fir@126837.6]
  wire [8:0] _GEN_3; // @[DMI.scala 112:64:chipyard.TestHarness.RocketConfig.fir@126837.6]
  wire [2:0] _GEN_7; // @[DMI.scala 112:64:chipyard.TestHarness.RocketConfig.fir@126837.6]
  wire  _T_102; // @[DMI.scala 121:53:chipyard.TestHarness.RocketConfig.fir@126861.4]
  assign addr = {io_dmi_req_bits_addr, 2'h0}; // @[DMI.scala 97:46:chipyard.TestHarness.RocketConfig.fir@126692.4]
  assign _T_100 = io_dmi_req_bits_op == 2'h2; // @[DMI.scala 111:30:chipyard.TestHarness.RocketConfig.fir@126824.4]
  assign _T_101 = io_dmi_req_bits_op == 2'h1; // @[DMI.scala 112:37:chipyard.TestHarness.RocketConfig.fir@126836.6]
  assign _GEN_2 = _T_101 ? 4'hf : 4'h0; // @[DMI.scala 112:64:chipyard.TestHarness.RocketConfig.fir@126837.6]
  assign _GEN_3 = _T_101 ? addr : 9'h40; // @[DMI.scala 112:64:chipyard.TestHarness.RocketConfig.fir@126837.6]
  assign _GEN_7 = _T_101 ? 3'h4 : 3'h1; // @[DMI.scala 112:64:chipyard.TestHarness.RocketConfig.fir@126837.6]
  assign _T_102 = auto_out_d_bits_corrupt | auto_out_d_bits_denied; // @[DMI.scala 121:53:chipyard.TestHarness.RocketConfig.fir@126861.4]
  assign auto_out_a_valid = io_dmi_req_valid; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@126689.4]
  assign auto_out_a_bits_opcode = _T_100 ? 3'h0 : _GEN_7; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@126689.4]
  assign auto_out_a_bits_address = _T_100 ? addr : _GEN_3; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@126689.4]
  assign auto_out_a_bits_mask = _T_100 ? 4'hf : _GEN_2; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@126689.4]
  assign auto_out_a_bits_data = _T_100 ? io_dmi_req_bits_data : 32'h0; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@126689.4]
  assign auto_out_d_ready = io_dmi_resp_ready; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@126689.4]
  assign io_dmi_req_ready = auto_out_a_ready; // @[DMI.scala 117:22:chipyard.TestHarness.RocketConfig.fir@126858.4]
  assign io_dmi_resp_valid = auto_out_d_valid; // @[DMI.scala 119:28:chipyard.TestHarness.RocketConfig.fir@126859.4]
  assign io_dmi_resp_bits_data = auto_out_d_bits_data; // @[DMI.scala 122:28:chipyard.TestHarness.RocketConfig.fir@126864.4]
  assign io_dmi_resp_bits_resp = {{1'd0}, _T_102}; // @[DMI.scala 121:28:chipyard.TestHarness.RocketConfig.fir@126863.4]
endmodule
