module ClockGroupAggregator( // @[:chipyard.TestHarness.RocketConfig.fir@43.2]
  input   auto_in_member_5_clock, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  input   auto_in_member_5_reset, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  input   auto_in_member_4_clock, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  input   auto_in_member_4_reset, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  input   auto_in_member_3_clock, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  input   auto_in_member_3_reset, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  input   auto_in_member_2_clock, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  input   auto_in_member_2_reset, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  input   auto_in_member_1_clock, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  input   auto_in_member_1_reset, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  input   auto_in_member_0_clock, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  input   auto_in_member_0_reset, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  output  auto_out_3_member_1_clock, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  output  auto_out_3_member_1_reset, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  output  auto_out_3_member_0_clock, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  output  auto_out_3_member_0_reset, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  output  auto_out_2_member_0_clock, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  output  auto_out_2_member_0_reset, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  output  auto_out_1_member_1_clock, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  output  auto_out_1_member_1_reset, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  output  auto_out_1_member_0_clock, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  output  auto_out_1_member_0_reset, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  output  auto_out_0_member_0_clock, // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
  output  auto_out_0_member_0_reset // @[:chipyard.TestHarness.RocketConfig.fir@44.4]
);
  assign auto_out_3_member_1_clock = auto_in_member_5_clock; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@67.4]
  assign auto_out_3_member_1_reset = auto_in_member_5_reset; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@67.4]
  assign auto_out_3_member_0_clock = auto_in_member_4_clock; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@67.4]
  assign auto_out_3_member_0_reset = auto_in_member_4_reset; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@67.4]
  assign auto_out_2_member_0_clock = auto_in_member_3_clock; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@66.4]
  assign auto_out_2_member_0_reset = auto_in_member_3_reset; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@66.4]
  assign auto_out_1_member_1_clock = auto_in_member_2_clock; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@65.4]
  assign auto_out_1_member_1_reset = auto_in_member_2_reset; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@65.4]
  assign auto_out_1_member_0_clock = auto_in_member_1_clock; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@65.4]
  assign auto_out_1_member_0_reset = auto_in_member_1_reset; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@65.4]
  assign auto_out_0_member_0_clock = auto_in_member_0_clock; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@64.4]
  assign auto_out_0_member_0_reset = auto_in_member_0_reset; // @[LazyModule.scala 181:49:chipyard.TestHarness.RocketConfig.fir@64.4]
endmodule
