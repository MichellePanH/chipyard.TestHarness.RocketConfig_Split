module ALU( // @[:chipyard.TestHarness.RocketConfig.fir@249564.2]
  input         io_dw, // @[:chipyard.TestHarness.RocketConfig.fir@249567.4]
  input  [3:0]  io_fn, // @[:chipyard.TestHarness.RocketConfig.fir@249567.4]
  input  [63:0] io_in2, // @[:chipyard.TestHarness.RocketConfig.fir@249567.4]
  input  [63:0] io_in1, // @[:chipyard.TestHarness.RocketConfig.fir@249567.4]
  output [63:0] io_out, // @[:chipyard.TestHarness.RocketConfig.fir@249567.4]
  output [63:0] io_adder_out, // @[:chipyard.TestHarness.RocketConfig.fir@249567.4]
  output        io_cmp_out // @[:chipyard.TestHarness.RocketConfig.fir@249567.4]
);
  wire [63:0] _T_1; // @[ALU.scala 62:35:chipyard.TestHarness.RocketConfig.fir@249573.4]
  wire [63:0] in2_inv; // @[ALU.scala 62:20:chipyard.TestHarness.RocketConfig.fir@249574.4]
  wire [63:0] in1_xor_in2; // @[ALU.scala 63:28:chipyard.TestHarness.RocketConfig.fir@249575.4]
  wire [63:0] _T_3; // @[ALU.scala 64:26:chipyard.TestHarness.RocketConfig.fir@249577.4]
  wire [63:0] _GEN_1; // @[ALU.scala 64:36:chipyard.TestHarness.RocketConfig.fir@249579.4]
  wire  _T_9; // @[ALU.scala 68:24:chipyard.TestHarness.RocketConfig.fir@249584.4]
  wire  _T_14; // @[ALU.scala 69:8:chipyard.TestHarness.RocketConfig.fir@249589.4]
  wire  slt; // @[ALU.scala 68:8:chipyard.TestHarness.RocketConfig.fir@249590.4]
  wire  _T_17; // @[ALU.scala 44:26:chipyard.TestHarness.RocketConfig.fir@249593.4]
  wire  _T_18; // @[ALU.scala 70:68:chipyard.TestHarness.RocketConfig.fir@249594.4]
  wire  _T_19; // @[ALU.scala 70:41:chipyard.TestHarness.RocketConfig.fir@249595.4]
  wire  _T_23; // @[ALU.scala 77:46:chipyard.TestHarness.RocketConfig.fir@249600.4]
  wire [31:0] _T_25; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@249602.4]
  wire [31:0] _T_28; // @[ALU.scala 78:24:chipyard.TestHarness.RocketConfig.fir@249605.4]
  wire  _T_31; // @[ALU.scala 79:33:chipyard.TestHarness.RocketConfig.fir@249608.4]
  wire [5:0] shamt; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@249610.4]
  wire [63:0] shin_r; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@249612.4]
  wire  _T_34; // @[ALU.scala 82:24:chipyard.TestHarness.RocketConfig.fir@249613.4]
  wire  _T_35; // @[ALU.scala 82:44:chipyard.TestHarness.RocketConfig.fir@249614.4]
  wire  _T_36; // @[ALU.scala 82:35:chipyard.TestHarness.RocketConfig.fir@249615.4]
  wire [63:0] _T_40; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249619.4]
  wire [63:0] _T_42; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249621.4]
  wire [63:0] _T_44; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249623.4]
  wire [63:0] _T_45; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249624.4]
  wire [63:0] _GEN_2; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249629.4]
  wire [63:0] _T_50; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249629.4]
  wire [63:0] _T_52; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249631.4]
  wire [63:0] _T_54; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249633.4]
  wire [63:0] _T_55; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249634.4]
  wire [63:0] _GEN_3; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249639.4]
  wire [63:0] _T_60; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249639.4]
  wire [63:0] _T_62; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249641.4]
  wire [63:0] _T_64; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249643.4]
  wire [63:0] _T_65; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249644.4]
  wire [63:0] _GEN_4; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249649.4]
  wire [63:0] _T_70; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249649.4]
  wire [63:0] _T_72; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249651.4]
  wire [63:0] _T_74; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249653.4]
  wire [63:0] _T_75; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249654.4]
  wire [63:0] _GEN_5; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249659.4]
  wire [63:0] _T_80; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249659.4]
  wire [63:0] _T_82; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249661.4]
  wire [63:0] _T_84; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249663.4]
  wire [63:0] _T_85; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249664.4]
  wire [63:0] _GEN_6; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249669.4]
  wire [63:0] _T_90; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249669.4]
  wire [63:0] _T_92; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249671.4]
  wire [63:0] _T_94; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249673.4]
  wire [63:0] _T_95; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249674.4]
  wire [63:0] shin; // @[ALU.scala 82:17:chipyard.TestHarness.RocketConfig.fir@249675.4]
  wire  _T_98; // @[ALU.scala 83:35:chipyard.TestHarness.RocketConfig.fir@249678.4]
  wire [64:0] _T_100; // @[ALU.scala 83:57:chipyard.TestHarness.RocketConfig.fir@249680.4]
  wire [64:0] _T_101; // @[ALU.scala 83:64:chipyard.TestHarness.RocketConfig.fir@249681.4]
  wire [63:0] shout_r; // @[ALU.scala 83:73:chipyard.TestHarness.RocketConfig.fir@249682.4]
  wire [63:0] _T_105; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249686.4]
  wire [63:0] _T_107; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249688.4]
  wire [63:0] _T_109; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249690.4]
  wire [63:0] _T_110; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249691.4]
  wire [63:0] _GEN_7; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249696.4]
  wire [63:0] _T_115; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249696.4]
  wire [63:0] _T_117; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249698.4]
  wire [63:0] _T_119; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249700.4]
  wire [63:0] _T_120; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249701.4]
  wire [63:0] _GEN_8; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249706.4]
  wire [63:0] _T_125; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249706.4]
  wire [63:0] _T_127; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249708.4]
  wire [63:0] _T_129; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249710.4]
  wire [63:0] _T_130; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249711.4]
  wire [63:0] _GEN_9; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249716.4]
  wire [63:0] _T_135; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249716.4]
  wire [63:0] _T_137; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249718.4]
  wire [63:0] _T_139; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249720.4]
  wire [63:0] _T_140; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249721.4]
  wire [63:0] _GEN_10; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249726.4]
  wire [63:0] _T_145; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249726.4]
  wire [63:0] _T_147; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249728.4]
  wire [63:0] _T_149; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249730.4]
  wire [63:0] _T_150; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249731.4]
  wire [63:0] _GEN_11; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249736.4]
  wire [63:0] _T_155; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249736.4]
  wire [63:0] _T_157; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249738.4]
  wire [63:0] _T_159; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249740.4]
  wire [63:0] shout_l; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249741.4]
  wire [63:0] _T_163; // @[ALU.scala 85:18:chipyard.TestHarness.RocketConfig.fir@249745.4]
  wire  _T_164; // @[ALU.scala 86:25:chipyard.TestHarness.RocketConfig.fir@249746.4]
  wire [63:0] _T_165; // @[ALU.scala 86:18:chipyard.TestHarness.RocketConfig.fir@249747.4]
  wire [63:0] shout; // @[ALU.scala 85:74:chipyard.TestHarness.RocketConfig.fir@249748.4]
  wire  _T_166; // @[ALU.scala 89:25:chipyard.TestHarness.RocketConfig.fir@249749.4]
  wire  _T_167; // @[ALU.scala 89:45:chipyard.TestHarness.RocketConfig.fir@249750.4]
  wire  _T_168; // @[ALU.scala 89:36:chipyard.TestHarness.RocketConfig.fir@249751.4]
  wire [63:0] _T_169; // @[ALU.scala 89:18:chipyard.TestHarness.RocketConfig.fir@249752.4]
  wire  _T_171; // @[ALU.scala 90:44:chipyard.TestHarness.RocketConfig.fir@249754.4]
  wire  _T_172; // @[ALU.scala 90:35:chipyard.TestHarness.RocketConfig.fir@249755.4]
  wire [63:0] _T_173; // @[ALU.scala 90:63:chipyard.TestHarness.RocketConfig.fir@249756.4]
  wire [63:0] _T_174; // @[ALU.scala 90:18:chipyard.TestHarness.RocketConfig.fir@249757.4]
  wire [63:0] logic_; // @[ALU.scala 89:78:chipyard.TestHarness.RocketConfig.fir@249758.4]
  wire  _T_175; // @[ALU.scala 41:30:chipyard.TestHarness.RocketConfig.fir@249759.4]
  wire  _T_176; // @[ALU.scala 91:35:chipyard.TestHarness.RocketConfig.fir@249760.4]
  wire [63:0] _GEN_12; // @[ALU.scala 91:43:chipyard.TestHarness.RocketConfig.fir@249761.4]
  wire [63:0] _T_177; // @[ALU.scala 91:43:chipyard.TestHarness.RocketConfig.fir@249761.4]
  wire [63:0] shift_logic; // @[ALU.scala 91:51:chipyard.TestHarness.RocketConfig.fir@249762.4]
  wire  _T_178; // @[ALU.scala 92:23:chipyard.TestHarness.RocketConfig.fir@249763.4]
  wire  _T_179; // @[ALU.scala 92:43:chipyard.TestHarness.RocketConfig.fir@249764.4]
  wire  _T_180; // @[ALU.scala 92:34:chipyard.TestHarness.RocketConfig.fir@249765.4]
  wire [63:0] out; // @[ALU.scala 92:16:chipyard.TestHarness.RocketConfig.fir@249766.4]
  wire  _T_181; // @[ALU.scala 97:17:chipyard.TestHarness.RocketConfig.fir@249768.4]
  wire [31:0] _T_184; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@249772.6]
  wire [63:0] _T_186; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@249774.6]
  assign _T_1 = ~io_in2; // @[ALU.scala 62:35:chipyard.TestHarness.RocketConfig.fir@249573.4]
  assign in2_inv = io_fn[3] ? _T_1 : io_in2; // @[ALU.scala 62:20:chipyard.TestHarness.RocketConfig.fir@249574.4]
  assign in1_xor_in2 = io_in1 ^ in2_inv; // @[ALU.scala 63:28:chipyard.TestHarness.RocketConfig.fir@249575.4]
  assign _T_3 = io_in1 + in2_inv; // @[ALU.scala 64:26:chipyard.TestHarness.RocketConfig.fir@249577.4]
  assign _GEN_1 = {{63'd0}, io_fn[3]}; // @[ALU.scala 64:36:chipyard.TestHarness.RocketConfig.fir@249579.4]
  assign _T_9 = io_in1[63] == io_in2[63]; // @[ALU.scala 68:24:chipyard.TestHarness.RocketConfig.fir@249584.4]
  assign _T_14 = io_fn[1] ? io_in2[63] : io_in1[63]; // @[ALU.scala 69:8:chipyard.TestHarness.RocketConfig.fir@249589.4]
  assign slt = _T_9 ? io_adder_out[63] : _T_14; // @[ALU.scala 68:8:chipyard.TestHarness.RocketConfig.fir@249590.4]
  assign _T_17 = ~io_fn[3]; // @[ALU.scala 44:26:chipyard.TestHarness.RocketConfig.fir@249593.4]
  assign _T_18 = in1_xor_in2 == 64'h0; // @[ALU.scala 70:68:chipyard.TestHarness.RocketConfig.fir@249594.4]
  assign _T_19 = _T_17 ? _T_18 : slt; // @[ALU.scala 70:41:chipyard.TestHarness.RocketConfig.fir@249595.4]
  assign _T_23 = io_fn[3] & io_in1[31]; // @[ALU.scala 77:46:chipyard.TestHarness.RocketConfig.fir@249600.4]
  assign _T_25 = _T_23 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@249602.4]
  assign _T_28 = io_dw ? io_in1[63:32] : _T_25; // @[ALU.scala 78:24:chipyard.TestHarness.RocketConfig.fir@249605.4]
  assign _T_31 = io_in2[5] & io_dw; // @[ALU.scala 79:33:chipyard.TestHarness.RocketConfig.fir@249608.4]
  assign shamt = {_T_31,io_in2[4:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@249610.4]
  assign shin_r = {_T_28,io_in1[31:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@249612.4]
  assign _T_34 = io_fn == 4'h5; // @[ALU.scala 82:24:chipyard.TestHarness.RocketConfig.fir@249613.4]
  assign _T_35 = io_fn == 4'hb; // @[ALU.scala 82:44:chipyard.TestHarness.RocketConfig.fir@249614.4]
  assign _T_36 = _T_34 | _T_35; // @[ALU.scala 82:35:chipyard.TestHarness.RocketConfig.fir@249615.4]
  assign _T_40 = {{32'd0}, shin_r[63:32]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249619.4]
  assign _T_42 = {shin_r[31:0], 32'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249621.4]
  assign _T_44 = _T_42 & 64'hffffffff00000000; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249623.4]
  assign _T_45 = _T_40 | _T_44; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249624.4]
  assign _GEN_2 = {{16'd0}, _T_45[63:16]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249629.4]
  assign _T_50 = _GEN_2 & 64'hffff0000ffff; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249629.4]
  assign _T_52 = {_T_45[47:0], 16'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249631.4]
  assign _T_54 = _T_52 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249633.4]
  assign _T_55 = _T_50 | _T_54; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249634.4]
  assign _GEN_3 = {{8'd0}, _T_55[63:8]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249639.4]
  assign _T_60 = _GEN_3 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249639.4]
  assign _T_62 = {_T_55[55:0], 8'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249641.4]
  assign _T_64 = _T_62 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249643.4]
  assign _T_65 = _T_60 | _T_64; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249644.4]
  assign _GEN_4 = {{4'd0}, _T_65[63:4]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249649.4]
  assign _T_70 = _GEN_4 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249649.4]
  assign _T_72 = {_T_65[59:0], 4'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249651.4]
  assign _T_74 = _T_72 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249653.4]
  assign _T_75 = _T_70 | _T_74; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249654.4]
  assign _GEN_5 = {{2'd0}, _T_75[63:2]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249659.4]
  assign _T_80 = _GEN_5 & 64'h3333333333333333; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249659.4]
  assign _T_82 = {_T_75[61:0], 2'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249661.4]
  assign _T_84 = _T_82 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249663.4]
  assign _T_85 = _T_80 | _T_84; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249664.4]
  assign _GEN_6 = {{1'd0}, _T_85[63:1]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249669.4]
  assign _T_90 = _GEN_6 & 64'h5555555555555555; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249669.4]
  assign _T_92 = {_T_85[62:0], 1'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249671.4]
  assign _T_94 = _T_92 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249673.4]
  assign _T_95 = _T_90 | _T_94; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249674.4]
  assign shin = _T_36 ? shin_r : _T_95; // @[ALU.scala 82:17:chipyard.TestHarness.RocketConfig.fir@249675.4]
  assign _T_98 = io_fn[3] & shin[63]; // @[ALU.scala 83:35:chipyard.TestHarness.RocketConfig.fir@249678.4]
  assign _T_100 = {_T_98,shin}; // @[ALU.scala 83:57:chipyard.TestHarness.RocketConfig.fir@249680.4]
  assign _T_101 = $signed(_T_100) >>> shamt; // @[ALU.scala 83:64:chipyard.TestHarness.RocketConfig.fir@249681.4]
  assign shout_r = _T_101[63:0]; // @[ALU.scala 83:73:chipyard.TestHarness.RocketConfig.fir@249682.4]
  assign _T_105 = {{32'd0}, shout_r[63:32]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249686.4]
  assign _T_107 = {shout_r[31:0], 32'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249688.4]
  assign _T_109 = _T_107 & 64'hffffffff00000000; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249690.4]
  assign _T_110 = _T_105 | _T_109; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249691.4]
  assign _GEN_7 = {{16'd0}, _T_110[63:16]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249696.4]
  assign _T_115 = _GEN_7 & 64'hffff0000ffff; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249696.4]
  assign _T_117 = {_T_110[47:0], 16'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249698.4]
  assign _T_119 = _T_117 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249700.4]
  assign _T_120 = _T_115 | _T_119; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249701.4]
  assign _GEN_8 = {{8'd0}, _T_120[63:8]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249706.4]
  assign _T_125 = _GEN_8 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249706.4]
  assign _T_127 = {_T_120[55:0], 8'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249708.4]
  assign _T_129 = _T_127 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249710.4]
  assign _T_130 = _T_125 | _T_129; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249711.4]
  assign _GEN_9 = {{4'd0}, _T_130[63:4]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249716.4]
  assign _T_135 = _GEN_9 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249716.4]
  assign _T_137 = {_T_130[59:0], 4'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249718.4]
  assign _T_139 = _T_137 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249720.4]
  assign _T_140 = _T_135 | _T_139; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249721.4]
  assign _GEN_10 = {{2'd0}, _T_140[63:2]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249726.4]
  assign _T_145 = _GEN_10 & 64'h3333333333333333; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249726.4]
  assign _T_147 = {_T_140[61:0], 2'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249728.4]
  assign _T_149 = _T_147 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249730.4]
  assign _T_150 = _T_145 | _T_149; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249731.4]
  assign _GEN_11 = {{1'd0}, _T_150[63:1]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249736.4]
  assign _T_155 = _GEN_11 & 64'h5555555555555555; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@249736.4]
  assign _T_157 = {_T_150[62:0], 1'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@249738.4]
  assign _T_159 = _T_157 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@249740.4]
  assign shout_l = _T_155 | _T_159; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@249741.4]
  assign _T_163 = _T_36 ? shout_r : 64'h0; // @[ALU.scala 85:18:chipyard.TestHarness.RocketConfig.fir@249745.4]
  assign _T_164 = io_fn == 4'h1; // @[ALU.scala 86:25:chipyard.TestHarness.RocketConfig.fir@249746.4]
  assign _T_165 = _T_164 ? shout_l : 64'h0; // @[ALU.scala 86:18:chipyard.TestHarness.RocketConfig.fir@249747.4]
  assign shout = _T_163 | _T_165; // @[ALU.scala 85:74:chipyard.TestHarness.RocketConfig.fir@249748.4]
  assign _T_166 = io_fn == 4'h4; // @[ALU.scala 89:25:chipyard.TestHarness.RocketConfig.fir@249749.4]
  assign _T_167 = io_fn == 4'h6; // @[ALU.scala 89:45:chipyard.TestHarness.RocketConfig.fir@249750.4]
  assign _T_168 = _T_166 | _T_167; // @[ALU.scala 89:36:chipyard.TestHarness.RocketConfig.fir@249751.4]
  assign _T_169 = _T_168 ? in1_xor_in2 : 64'h0; // @[ALU.scala 89:18:chipyard.TestHarness.RocketConfig.fir@249752.4]
  assign _T_171 = io_fn == 4'h7; // @[ALU.scala 90:44:chipyard.TestHarness.RocketConfig.fir@249754.4]
  assign _T_172 = _T_167 | _T_171; // @[ALU.scala 90:35:chipyard.TestHarness.RocketConfig.fir@249755.4]
  assign _T_173 = io_in1 & io_in2; // @[ALU.scala 90:63:chipyard.TestHarness.RocketConfig.fir@249756.4]
  assign _T_174 = _T_172 ? _T_173 : 64'h0; // @[ALU.scala 90:18:chipyard.TestHarness.RocketConfig.fir@249757.4]
  assign logic_ = _T_169 | _T_174; // @[ALU.scala 89:78:chipyard.TestHarness.RocketConfig.fir@249758.4]
  assign _T_175 = io_fn >= 4'hc; // @[ALU.scala 41:30:chipyard.TestHarness.RocketConfig.fir@249759.4]
  assign _T_176 = _T_175 & slt; // @[ALU.scala 91:35:chipyard.TestHarness.RocketConfig.fir@249760.4]
  assign _GEN_12 = {{63'd0}, _T_176}; // @[ALU.scala 91:43:chipyard.TestHarness.RocketConfig.fir@249761.4]
  assign _T_177 = _GEN_12 | logic_; // @[ALU.scala 91:43:chipyard.TestHarness.RocketConfig.fir@249761.4]
  assign shift_logic = _T_177 | shout; // @[ALU.scala 91:51:chipyard.TestHarness.RocketConfig.fir@249762.4]
  assign _T_178 = io_fn == 4'h0; // @[ALU.scala 92:23:chipyard.TestHarness.RocketConfig.fir@249763.4]
  assign _T_179 = io_fn == 4'ha; // @[ALU.scala 92:43:chipyard.TestHarness.RocketConfig.fir@249764.4]
  assign _T_180 = _T_178 | _T_179; // @[ALU.scala 92:34:chipyard.TestHarness.RocketConfig.fir@249765.4]
  assign out = _T_180 ? io_adder_out : shift_logic; // @[ALU.scala 92:16:chipyard.TestHarness.RocketConfig.fir@249766.4]
  assign _T_181 = ~io_dw; // @[ALU.scala 97:17:chipyard.TestHarness.RocketConfig.fir@249768.4]
  assign _T_184 = out[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@249772.6]
  assign _T_186 = {_T_184,out[31:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@249774.6]
  assign io_out = _T_181 ? _T_186 : out; // @[ALU.scala 94:10:chipyard.TestHarness.RocketConfig.fir@249767.4 ALU.scala 97:37:chipyard.TestHarness.RocketConfig.fir@249775.6]
  assign io_adder_out = _T_3 + _GEN_1; // @[ALU.scala 64:16:chipyard.TestHarness.RocketConfig.fir@249581.4]
  assign io_cmp_out = io_fn[0] ^ _T_19; // @[ALU.scala 70:14:chipyard.TestHarness.RocketConfig.fir@249597.4]
endmodule
