module package_Anon_118( // @[:chipyard.TestHarness.RocketConfig.fir@240856.2]
  input  [53:0] io_x_ppn, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  input         io_x_d, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  input         io_x_a, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  input         io_x_g, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  input         io_x_u, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  input         io_x_x, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  input         io_x_w, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  input         io_x_r, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  input         io_x_v, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  output [53:0] io_y_ppn, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  output        io_y_d, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  output        io_y_a, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  output        io_y_g, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  output        io_y_u, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  output        io_y_x, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  output        io_y_w, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  output        io_y_r, // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
  output        io_y_v // @[:chipyard.TestHarness.RocketConfig.fir@240859.4]
);
  assign io_y_ppn = io_x_ppn; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@240864.4]
  assign io_y_d = io_x_d; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@240864.4]
  assign io_y_a = io_x_a; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@240864.4]
  assign io_y_g = io_x_g; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@240864.4]
  assign io_y_u = io_x_u; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@240864.4]
  assign io_y_x = io_x_x; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@240864.4]
  assign io_y_w = io_x_w; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@240864.4]
  assign io_y_r = io_x_r; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@240864.4]
  assign io_y_v = io_x_v; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@240864.4]
endmodule
