module PMPChecker_2( // @[:chipyard.TestHarness.RocketConfig.fir@219627.2]
  input  [1:0]  io_prv, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_0_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [1:0]  io_pmp_0_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_0_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_0_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_0_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [29:0] io_pmp_0_addr, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [31:0] io_pmp_0_mask, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_1_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [1:0]  io_pmp_1_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_1_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_1_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_1_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [29:0] io_pmp_1_addr, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [31:0] io_pmp_1_mask, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_2_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [1:0]  io_pmp_2_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_2_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_2_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_2_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [29:0] io_pmp_2_addr, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [31:0] io_pmp_2_mask, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_3_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [1:0]  io_pmp_3_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_3_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_3_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_3_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [29:0] io_pmp_3_addr, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [31:0] io_pmp_3_mask, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_4_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [1:0]  io_pmp_4_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_4_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_4_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_4_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [29:0] io_pmp_4_addr, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [31:0] io_pmp_4_mask, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_5_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [1:0]  io_pmp_5_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_5_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_5_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_5_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [29:0] io_pmp_5_addr, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [31:0] io_pmp_5_mask, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_6_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [1:0]  io_pmp_6_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_6_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_6_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_6_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [29:0] io_pmp_6_addr, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [31:0] io_pmp_6_mask, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_7_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [1:0]  io_pmp_7_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_7_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_7_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input         io_pmp_7_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [29:0] io_pmp_7_addr, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [31:0] io_pmp_7_mask, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  input  [31:0] io_addr, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  output        io_r, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  output        io_w, // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
  output        io_x // @[:chipyard.TestHarness.RocketConfig.fir@219630.4]
);
  wire  default_; // @[PMP.scala 157:56:chipyard.TestHarness.RocketConfig.fir@219632.4]
  wire [31:0] _T_2; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@219655.4]
  wire [31:0] _T_3; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@219656.4]
  wire [31:0] _T_4; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@219657.4]
  wire [31:0] _T_5; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@219658.4]
  wire [31:0] _T_6; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@219659.4]
  wire [31:0] _T_7; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@219660.4]
  wire [31:0] _T_8; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@219661.4]
  wire  _T_9; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@219662.4]
  wire [31:0] _T_15; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@219668.4]
  wire [31:0] _T_16; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@219669.4]
  wire [31:0] _T_17; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@219670.4]
  wire [31:0] _T_18; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@219671.4]
  wire  _T_19; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@219672.4]
  wire  _T_20; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@219673.4]
  wire  _T_25; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@219678.4]
  wire  _T_26; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@219679.4]
  wire  _T_27; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@219680.4]
  wire  _T_28; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@219681.4]
  wire  _T_29; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@219682.4]
  wire  _T_30; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@219683.4]
  wire  _T_82; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@219743.4]
  wire  _T_84; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@219746.4]
  wire  _T_86; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@219749.4]
  wire  _T_88_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219752.4]
  wire  _T_88_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219752.4]
  wire  _T_88_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219752.4]
  wire [31:0] _T_94; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@219758.4]
  wire [31:0] _T_95; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@219759.4]
  wire [31:0] _T_96; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@219760.4]
  wire  _T_97; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@219761.4]
  wire [31:0] _T_103; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@219767.4]
  wire [31:0] _T_104; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@219768.4]
  wire [31:0] _T_105; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@219769.4]
  wire [31:0] _T_106; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@219770.4]
  wire  _T_107; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@219771.4]
  wire  _T_108; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@219772.4]
  wire  _T_114; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@219778.4]
  wire  _T_115; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@219779.4]
  wire  _T_116; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@219780.4]
  wire  _T_117; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@219781.4]
  wire  _T_118; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@219782.4]
  wire  _T_170; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@219842.4]
  wire  _T_172; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@219845.4]
  wire  _T_174; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@219848.4]
  wire  _T_176_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219851.4]
  wire  _T_176_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219851.4]
  wire  _T_176_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219851.4]
  wire [31:0] _T_182; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@219857.4]
  wire [31:0] _T_183; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@219858.4]
  wire [31:0] _T_184; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@219859.4]
  wire  _T_185; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@219860.4]
  wire [31:0] _T_191; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@219866.4]
  wire [31:0] _T_192; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@219867.4]
  wire [31:0] _T_193; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@219868.4]
  wire [31:0] _T_194; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@219869.4]
  wire  _T_195; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@219870.4]
  wire  _T_196; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@219871.4]
  wire  _T_202; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@219877.4]
  wire  _T_203; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@219878.4]
  wire  _T_204; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@219879.4]
  wire  _T_205; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@219880.4]
  wire  _T_206; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@219881.4]
  wire  _T_258; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@219941.4]
  wire  _T_260; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@219944.4]
  wire  _T_262; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@219947.4]
  wire  _T_264_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219950.4]
  wire  _T_264_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219950.4]
  wire  _T_264_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219950.4]
  wire [31:0] _T_270; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@219956.4]
  wire [31:0] _T_271; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@219957.4]
  wire [31:0] _T_272; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@219958.4]
  wire  _T_273; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@219959.4]
  wire [31:0] _T_279; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@219965.4]
  wire [31:0] _T_280; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@219966.4]
  wire [31:0] _T_281; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@219967.4]
  wire [31:0] _T_282; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@219968.4]
  wire  _T_283; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@219969.4]
  wire  _T_284; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@219970.4]
  wire  _T_290; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@219976.4]
  wire  _T_291; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@219977.4]
  wire  _T_292; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@219978.4]
  wire  _T_293; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@219979.4]
  wire  _T_294; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@219980.4]
  wire  _T_346; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@220040.4]
  wire  _T_348; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@220043.4]
  wire  _T_350; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@220046.4]
  wire  _T_352_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220049.4]
  wire  _T_352_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220049.4]
  wire  _T_352_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220049.4]
  wire [31:0] _T_358; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@220055.4]
  wire [31:0] _T_359; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@220056.4]
  wire [31:0] _T_360; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@220057.4]
  wire  _T_361; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@220058.4]
  wire [31:0] _T_367; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@220064.4]
  wire [31:0] _T_368; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@220065.4]
  wire [31:0] _T_369; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@220066.4]
  wire [31:0] _T_370; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@220067.4]
  wire  _T_371; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@220068.4]
  wire  _T_372; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@220069.4]
  wire  _T_378; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@220075.4]
  wire  _T_379; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@220076.4]
  wire  _T_380; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@220077.4]
  wire  _T_381; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@220078.4]
  wire  _T_382; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@220079.4]
  wire  _T_434; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@220139.4]
  wire  _T_436; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@220142.4]
  wire  _T_438; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@220145.4]
  wire  _T_440_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220148.4]
  wire  _T_440_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220148.4]
  wire  _T_440_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220148.4]
  wire [31:0] _T_446; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@220154.4]
  wire [31:0] _T_447; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@220155.4]
  wire [31:0] _T_448; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@220156.4]
  wire  _T_449; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@220157.4]
  wire [31:0] _T_455; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@220163.4]
  wire [31:0] _T_456; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@220164.4]
  wire [31:0] _T_457; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@220165.4]
  wire [31:0] _T_458; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@220166.4]
  wire  _T_459; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@220167.4]
  wire  _T_460; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@220168.4]
  wire  _T_466; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@220174.4]
  wire  _T_467; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@220175.4]
  wire  _T_468; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@220176.4]
  wire  _T_469; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@220177.4]
  wire  _T_470; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@220178.4]
  wire  _T_522; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@220238.4]
  wire  _T_524; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@220241.4]
  wire  _T_526; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@220244.4]
  wire  _T_528_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220247.4]
  wire  _T_528_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220247.4]
  wire  _T_528_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220247.4]
  wire [31:0] _T_534; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@220253.4]
  wire [31:0] _T_535; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@220254.4]
  wire [31:0] _T_536; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@220255.4]
  wire  _T_537; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@220256.4]
  wire [31:0] _T_543; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@220262.4]
  wire [31:0] _T_544; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@220263.4]
  wire [31:0] _T_545; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@220264.4]
  wire [31:0] _T_546; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@220265.4]
  wire  _T_547; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@220266.4]
  wire  _T_548; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@220267.4]
  wire  _T_554; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@220273.4]
  wire  _T_555; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@220274.4]
  wire  _T_556; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@220275.4]
  wire  _T_557; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@220276.4]
  wire  _T_558; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@220277.4]
  wire  _T_610; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@220337.4]
  wire  _T_612; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@220340.4]
  wire  _T_614; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@220343.4]
  wire  _T_616_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220346.4]
  wire  _T_616_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220346.4]
  wire  _T_616_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220346.4]
  wire [31:0] _T_622; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@220352.4]
  wire [31:0] _T_623; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@220353.4]
  wire [31:0] _T_624; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@220354.4]
  wire  _T_625; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@220355.4]
  wire  _T_643; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@220373.4]
  wire  _T_644; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@220374.4]
  wire  _T_645; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@220375.4]
  wire  _T_646; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@220376.4]
  wire  _T_698; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@220436.4]
  wire  _T_700; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@220439.4]
  wire  _T_702; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@220442.4]
  assign default_ = io_prv > 2'h1; // @[PMP.scala 157:56:chipyard.TestHarness.RocketConfig.fir@219632.4]
  assign _T_2 = {io_pmp_7_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@219655.4]
  assign _T_3 = ~_T_2; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@219656.4]
  assign _T_4 = _T_3 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@219657.4]
  assign _T_5 = ~_T_4; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@219658.4]
  assign _T_6 = io_addr ^ _T_5; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@219659.4]
  assign _T_7 = ~io_pmp_7_mask; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@219660.4]
  assign _T_8 = _T_6 & _T_7; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@219661.4]
  assign _T_9 = _T_8 == 32'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@219662.4]
  assign _T_15 = {io_pmp_6_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@219668.4]
  assign _T_16 = ~_T_15; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@219669.4]
  assign _T_17 = _T_16 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@219670.4]
  assign _T_18 = ~_T_17; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@219671.4]
  assign _T_19 = io_addr < _T_18; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@219672.4]
  assign _T_20 = ~_T_19; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@219673.4]
  assign _T_25 = io_addr < _T_5; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@219678.4]
  assign _T_26 = _T_20 & _T_25; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@219679.4]
  assign _T_27 = io_pmp_7_cfg_a[0] & _T_26; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@219680.4]
  assign _T_28 = io_pmp_7_cfg_a[1] ? _T_9 : _T_27; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@219681.4]
  assign _T_29 = ~io_pmp_7_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@219682.4]
  assign _T_30 = default_ & _T_29; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@219683.4]
  assign _T_82 = io_pmp_7_cfg_r | _T_30; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@219743.4]
  assign _T_84 = io_pmp_7_cfg_w | _T_30; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@219746.4]
  assign _T_86 = io_pmp_7_cfg_x | _T_30; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@219749.4]
  assign _T_88_cfg_x = _T_28 ? _T_86 : default_; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219752.4]
  assign _T_88_cfg_w = _T_28 ? _T_84 : default_; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219752.4]
  assign _T_88_cfg_r = _T_28 ? _T_82 : default_; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219752.4]
  assign _T_94 = io_addr ^ _T_18; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@219758.4]
  assign _T_95 = ~io_pmp_6_mask; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@219759.4]
  assign _T_96 = _T_94 & _T_95; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@219760.4]
  assign _T_97 = _T_96 == 32'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@219761.4]
  assign _T_103 = {io_pmp_5_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@219767.4]
  assign _T_104 = ~_T_103; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@219768.4]
  assign _T_105 = _T_104 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@219769.4]
  assign _T_106 = ~_T_105; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@219770.4]
  assign _T_107 = io_addr < _T_106; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@219771.4]
  assign _T_108 = ~_T_107; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@219772.4]
  assign _T_114 = _T_108 & _T_19; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@219778.4]
  assign _T_115 = io_pmp_6_cfg_a[0] & _T_114; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@219779.4]
  assign _T_116 = io_pmp_6_cfg_a[1] ? _T_97 : _T_115; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@219780.4]
  assign _T_117 = ~io_pmp_6_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@219781.4]
  assign _T_118 = default_ & _T_117; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@219782.4]
  assign _T_170 = io_pmp_6_cfg_r | _T_118; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@219842.4]
  assign _T_172 = io_pmp_6_cfg_w | _T_118; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@219845.4]
  assign _T_174 = io_pmp_6_cfg_x | _T_118; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@219848.4]
  assign _T_176_cfg_x = _T_116 ? _T_174 : _T_88_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219851.4]
  assign _T_176_cfg_w = _T_116 ? _T_172 : _T_88_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219851.4]
  assign _T_176_cfg_r = _T_116 ? _T_170 : _T_88_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219851.4]
  assign _T_182 = io_addr ^ _T_106; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@219857.4]
  assign _T_183 = ~io_pmp_5_mask; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@219858.4]
  assign _T_184 = _T_182 & _T_183; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@219859.4]
  assign _T_185 = _T_184 == 32'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@219860.4]
  assign _T_191 = {io_pmp_4_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@219866.4]
  assign _T_192 = ~_T_191; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@219867.4]
  assign _T_193 = _T_192 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@219868.4]
  assign _T_194 = ~_T_193; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@219869.4]
  assign _T_195 = io_addr < _T_194; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@219870.4]
  assign _T_196 = ~_T_195; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@219871.4]
  assign _T_202 = _T_196 & _T_107; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@219877.4]
  assign _T_203 = io_pmp_5_cfg_a[0] & _T_202; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@219878.4]
  assign _T_204 = io_pmp_5_cfg_a[1] ? _T_185 : _T_203; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@219879.4]
  assign _T_205 = ~io_pmp_5_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@219880.4]
  assign _T_206 = default_ & _T_205; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@219881.4]
  assign _T_258 = io_pmp_5_cfg_r | _T_206; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@219941.4]
  assign _T_260 = io_pmp_5_cfg_w | _T_206; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@219944.4]
  assign _T_262 = io_pmp_5_cfg_x | _T_206; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@219947.4]
  assign _T_264_cfg_x = _T_204 ? _T_262 : _T_176_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219950.4]
  assign _T_264_cfg_w = _T_204 ? _T_260 : _T_176_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219950.4]
  assign _T_264_cfg_r = _T_204 ? _T_258 : _T_176_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@219950.4]
  assign _T_270 = io_addr ^ _T_194; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@219956.4]
  assign _T_271 = ~io_pmp_4_mask; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@219957.4]
  assign _T_272 = _T_270 & _T_271; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@219958.4]
  assign _T_273 = _T_272 == 32'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@219959.4]
  assign _T_279 = {io_pmp_3_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@219965.4]
  assign _T_280 = ~_T_279; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@219966.4]
  assign _T_281 = _T_280 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@219967.4]
  assign _T_282 = ~_T_281; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@219968.4]
  assign _T_283 = io_addr < _T_282; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@219969.4]
  assign _T_284 = ~_T_283; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@219970.4]
  assign _T_290 = _T_284 & _T_195; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@219976.4]
  assign _T_291 = io_pmp_4_cfg_a[0] & _T_290; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@219977.4]
  assign _T_292 = io_pmp_4_cfg_a[1] ? _T_273 : _T_291; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@219978.4]
  assign _T_293 = ~io_pmp_4_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@219979.4]
  assign _T_294 = default_ & _T_293; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@219980.4]
  assign _T_346 = io_pmp_4_cfg_r | _T_294; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@220040.4]
  assign _T_348 = io_pmp_4_cfg_w | _T_294; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@220043.4]
  assign _T_350 = io_pmp_4_cfg_x | _T_294; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@220046.4]
  assign _T_352_cfg_x = _T_292 ? _T_350 : _T_264_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220049.4]
  assign _T_352_cfg_w = _T_292 ? _T_348 : _T_264_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220049.4]
  assign _T_352_cfg_r = _T_292 ? _T_346 : _T_264_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220049.4]
  assign _T_358 = io_addr ^ _T_282; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@220055.4]
  assign _T_359 = ~io_pmp_3_mask; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@220056.4]
  assign _T_360 = _T_358 & _T_359; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@220057.4]
  assign _T_361 = _T_360 == 32'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@220058.4]
  assign _T_367 = {io_pmp_2_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@220064.4]
  assign _T_368 = ~_T_367; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@220065.4]
  assign _T_369 = _T_368 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@220066.4]
  assign _T_370 = ~_T_369; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@220067.4]
  assign _T_371 = io_addr < _T_370; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@220068.4]
  assign _T_372 = ~_T_371; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@220069.4]
  assign _T_378 = _T_372 & _T_283; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@220075.4]
  assign _T_379 = io_pmp_3_cfg_a[0] & _T_378; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@220076.4]
  assign _T_380 = io_pmp_3_cfg_a[1] ? _T_361 : _T_379; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@220077.4]
  assign _T_381 = ~io_pmp_3_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@220078.4]
  assign _T_382 = default_ & _T_381; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@220079.4]
  assign _T_434 = io_pmp_3_cfg_r | _T_382; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@220139.4]
  assign _T_436 = io_pmp_3_cfg_w | _T_382; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@220142.4]
  assign _T_438 = io_pmp_3_cfg_x | _T_382; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@220145.4]
  assign _T_440_cfg_x = _T_380 ? _T_438 : _T_352_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220148.4]
  assign _T_440_cfg_w = _T_380 ? _T_436 : _T_352_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220148.4]
  assign _T_440_cfg_r = _T_380 ? _T_434 : _T_352_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220148.4]
  assign _T_446 = io_addr ^ _T_370; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@220154.4]
  assign _T_447 = ~io_pmp_2_mask; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@220155.4]
  assign _T_448 = _T_446 & _T_447; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@220156.4]
  assign _T_449 = _T_448 == 32'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@220157.4]
  assign _T_455 = {io_pmp_1_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@220163.4]
  assign _T_456 = ~_T_455; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@220164.4]
  assign _T_457 = _T_456 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@220165.4]
  assign _T_458 = ~_T_457; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@220166.4]
  assign _T_459 = io_addr < _T_458; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@220167.4]
  assign _T_460 = ~_T_459; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@220168.4]
  assign _T_466 = _T_460 & _T_371; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@220174.4]
  assign _T_467 = io_pmp_2_cfg_a[0] & _T_466; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@220175.4]
  assign _T_468 = io_pmp_2_cfg_a[1] ? _T_449 : _T_467; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@220176.4]
  assign _T_469 = ~io_pmp_2_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@220177.4]
  assign _T_470 = default_ & _T_469; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@220178.4]
  assign _T_522 = io_pmp_2_cfg_r | _T_470; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@220238.4]
  assign _T_524 = io_pmp_2_cfg_w | _T_470; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@220241.4]
  assign _T_526 = io_pmp_2_cfg_x | _T_470; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@220244.4]
  assign _T_528_cfg_x = _T_468 ? _T_526 : _T_440_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220247.4]
  assign _T_528_cfg_w = _T_468 ? _T_524 : _T_440_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220247.4]
  assign _T_528_cfg_r = _T_468 ? _T_522 : _T_440_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220247.4]
  assign _T_534 = io_addr ^ _T_458; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@220253.4]
  assign _T_535 = ~io_pmp_1_mask; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@220254.4]
  assign _T_536 = _T_534 & _T_535; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@220255.4]
  assign _T_537 = _T_536 == 32'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@220256.4]
  assign _T_543 = {io_pmp_0_addr, 2'h0}; // @[PMP.scala 62:36:chipyard.TestHarness.RocketConfig.fir@220262.4]
  assign _T_544 = ~_T_543; // @[PMP.scala 62:29:chipyard.TestHarness.RocketConfig.fir@220263.4]
  assign _T_545 = _T_544 | 32'h3; // @[PMP.scala 62:48:chipyard.TestHarness.RocketConfig.fir@220264.4]
  assign _T_546 = ~_T_545; // @[PMP.scala 62:27:chipyard.TestHarness.RocketConfig.fir@220265.4]
  assign _T_547 = io_addr < _T_546; // @[PMP.scala 79:9:chipyard.TestHarness.RocketConfig.fir@220266.4]
  assign _T_548 = ~_T_547; // @[PMP.scala 90:5:chipyard.TestHarness.RocketConfig.fir@220267.4]
  assign _T_554 = _T_548 & _T_459; // @[PMP.scala 96:48:chipyard.TestHarness.RocketConfig.fir@220273.4]
  assign _T_555 = io_pmp_1_cfg_a[0] & _T_554; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@220274.4]
  assign _T_556 = io_pmp_1_cfg_a[1] ? _T_537 : _T_555; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@220275.4]
  assign _T_557 = ~io_pmp_1_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@220276.4]
  assign _T_558 = default_ & _T_557; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@220277.4]
  assign _T_610 = io_pmp_1_cfg_r | _T_558; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@220337.4]
  assign _T_612 = io_pmp_1_cfg_w | _T_558; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@220340.4]
  assign _T_614 = io_pmp_1_cfg_x | _T_558; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@220343.4]
  assign _T_616_cfg_x = _T_556 ? _T_614 : _T_528_cfg_x; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220346.4]
  assign _T_616_cfg_w = _T_556 ? _T_612 : _T_528_cfg_w; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220346.4]
  assign _T_616_cfg_r = _T_556 ? _T_610 : _T_528_cfg_r; // @[PMP.scala 186:8:chipyard.TestHarness.RocketConfig.fir@220346.4]
  assign _T_622 = io_addr ^ _T_546; // @[PMP.scala 65:47:chipyard.TestHarness.RocketConfig.fir@220352.4]
  assign _T_623 = ~io_pmp_0_mask; // @[PMP.scala 65:54:chipyard.TestHarness.RocketConfig.fir@220353.4]
  assign _T_624 = _T_622 & _T_623; // @[PMP.scala 65:52:chipyard.TestHarness.RocketConfig.fir@220354.4]
  assign _T_625 = _T_624 == 32'h0; // @[PMP.scala 65:58:chipyard.TestHarness.RocketConfig.fir@220355.4]
  assign _T_643 = io_pmp_0_cfg_a[0] & _T_547; // @[PMP.scala 134:61:chipyard.TestHarness.RocketConfig.fir@220373.4]
  assign _T_644 = io_pmp_0_cfg_a[1] ? _T_625 : _T_643; // @[PMP.scala 134:8:chipyard.TestHarness.RocketConfig.fir@220374.4]
  assign _T_645 = ~io_pmp_0_cfg_l; // @[PMP.scala 165:29:chipyard.TestHarness.RocketConfig.fir@220375.4]
  assign _T_646 = default_ & _T_645; // @[PMP.scala 165:26:chipyard.TestHarness.RocketConfig.fir@220376.4]
  assign _T_698 = io_pmp_0_cfg_r | _T_646; // @[PMP.scala 183:40:chipyard.TestHarness.RocketConfig.fir@220436.4]
  assign _T_700 = io_pmp_0_cfg_w | _T_646; // @[PMP.scala 184:40:chipyard.TestHarness.RocketConfig.fir@220439.4]
  assign _T_702 = io_pmp_0_cfg_x | _T_646; // @[PMP.scala 185:40:chipyard.TestHarness.RocketConfig.fir@220442.4]
  assign io_r = _T_644 ? _T_698 : _T_616_cfg_r; // @[PMP.scala 189:8:chipyard.TestHarness.RocketConfig.fir@220446.4]
  assign io_w = _T_644 ? _T_700 : _T_616_cfg_w; // @[PMP.scala 190:8:chipyard.TestHarness.RocketConfig.fir@220447.4]
  assign io_x = _T_644 ? _T_702 : _T_616_cfg_x; // @[PMP.scala 191:8:chipyard.TestHarness.RocketConfig.fir@220448.4]
endmodule
