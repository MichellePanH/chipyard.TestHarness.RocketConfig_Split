module RVCExpander( // @[:chipyard.TestHarness.RocketConfig.fir@242309.2]
  input  [31:0] io_in, // @[:chipyard.TestHarness.RocketConfig.fir@242312.4]
  output [31:0] io_out_bits, // @[:chipyard.TestHarness.RocketConfig.fir@242312.4]
  output [4:0]  io_out_rd, // @[:chipyard.TestHarness.RocketConfig.fir@242312.4]
  output [4:0]  io_out_rs1, // @[:chipyard.TestHarness.RocketConfig.fir@242312.4]
  output [4:0]  io_out_rs2, // @[:chipyard.TestHarness.RocketConfig.fir@242312.4]
  output [4:0]  io_out_rs3, // @[:chipyard.TestHarness.RocketConfig.fir@242312.4]
  output        io_rvc // @[:chipyard.TestHarness.RocketConfig.fir@242312.4]
);
  wire  _T_3; // @[RVC.scala 54:29:chipyard.TestHarness.RocketConfig.fir@242318.4]
  wire [6:0] _T_4; // @[RVC.scala 54:20:chipyard.TestHarness.RocketConfig.fir@242319.4]
  wire [4:0] _T_14; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242329.4]
  wire [29:0] _T_18; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242333.4]
  wire [7:0] _T_28; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242348.4]
  wire [4:0] _T_30; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242350.4]
  wire [27:0] _T_36; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242356.4]
  wire [6:0] _T_50; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242375.4]
  wire [26:0] _T_58; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242383.4]
  wire [27:0] _T_78; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242408.4]
  wire [26:0] _T_109; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242444.4]
  wire [27:0] _T_136; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242476.4]
  wire [26:0] _T_167; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242512.4]
  wire [27:0] _T_194; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242544.4]
  wire [6:0] _T_205; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@242560.4]
  wire [11:0] _T_207; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242562.4]
  wire [31:0] _T_213; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242568.4]
  wire  _T_221; // @[RVC.scala 78:24:chipyard.TestHarness.RocketConfig.fir@242581.4]
  wire [6:0] _T_222; // @[RVC.scala 78:20:chipyard.TestHarness.RocketConfig.fir@242582.4]
  wire [31:0] _T_233; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242593.4]
  wire [31:0] _T_249; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242614.4]
  wire  _T_260; // @[RVC.scala 91:29:chipyard.TestHarness.RocketConfig.fir@242630.4]
  wire [6:0] _T_261; // @[RVC.scala 91:20:chipyard.TestHarness.RocketConfig.fir@242631.4]
  wire [14:0] _T_264; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@242634.4]
  wire [31:0] _T_267; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242637.4]
  wire [31:0] _T_271; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242641.4]
  wire  _T_279; // @[RVC.scala 93:14:chipyard.TestHarness.RocketConfig.fir@242654.4]
  wire  _T_281; // @[RVC.scala 93:27:chipyard.TestHarness.RocketConfig.fir@242656.4]
  wire  _T_282; // @[RVC.scala 93:21:chipyard.TestHarness.RocketConfig.fir@242657.4]
  wire [6:0] _T_289; // @[RVC.scala 87:20:chipyard.TestHarness.RocketConfig.fir@242664.4]
  wire [2:0] _T_292; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@242667.4]
  wire [31:0] _T_307; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242682.4]
  wire [31:0] _T_314_bits; // @[RVC.scala 93:10:chipyard.TestHarness.RocketConfig.fir@242694.4]
  wire [4:0] _T_314_rd; // @[RVC.scala 93:10:chipyard.TestHarness.RocketConfig.fir@242694.4]
  wire [4:0] _T_314_rs2; // @[RVC.scala 93:10:chipyard.TestHarness.RocketConfig.fir@242694.4]
  wire [4:0] _T_314_rs3; // @[RVC.scala 93:10:chipyard.TestHarness.RocketConfig.fir@242694.4]
  wire [25:0] _T_325; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242705.4]
  wire [30:0] _GEN_0; // @[RVC.scala 100:23:chipyard.TestHarness.RocketConfig.fir@242717.4]
  wire [30:0] _T_337; // @[RVC.scala 100:23:chipyard.TestHarness.RocketConfig.fir@242717.4]
  wire [31:0] _T_350; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242730.4]
  wire [2:0] _T_353; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242733.4]
  wire  _T_354; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242734.4]
  wire [2:0] _T_355; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242735.4]
  wire  _T_356; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242736.4]
  wire [2:0] _T_357; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242737.4]
  wire  _T_358; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242738.4]
  wire [2:0] _T_359; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242739.4]
  wire  _T_360; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242740.4]
  wire [2:0] _T_361; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242741.4]
  wire  _T_362; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242742.4]
  wire [2:0] _T_363; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242743.4]
  wire  _T_364; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242744.4]
  wire [2:0] _T_365; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242745.4]
  wire  _T_366; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242746.4]
  wire [2:0] _T_367; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242747.4]
  wire  _T_369; // @[RVC.scala 104:30:chipyard.TestHarness.RocketConfig.fir@242749.4]
  wire [30:0] _T_370; // @[RVC.scala 104:22:chipyard.TestHarness.RocketConfig.fir@242750.4]
  wire [6:0] _T_372; // @[RVC.scala 105:22:chipyard.TestHarness.RocketConfig.fir@242752.4]
  wire [24:0] _T_382; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242762.4]
  wire [30:0] _GEN_1; // @[RVC.scala 106:43:chipyard.TestHarness.RocketConfig.fir@242763.4]
  wire [30:0] _T_383; // @[RVC.scala 106:43:chipyard.TestHarness.RocketConfig.fir@242763.4]
  wire  _T_385; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242765.4]
  wire [30:0] _T_386; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242766.4]
  wire  _T_387; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242767.4]
  wire [31:0] _T_388; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242768.4]
  wire  _T_389; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242769.4]
  wire [31:0] _T_390; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242770.4]
  wire [9:0] _T_401; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@242786.4]
  wire [20:0] _T_416; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242801.4]
  wire [31:0] _T_479; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242864.4]
  wire [4:0] _T_488; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@242878.4]
  wire [12:0] _T_497; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242887.4]
  wire [31:0] _T_546; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242936.4]
  wire [31:0] _T_613; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243008.4]
  wire [6:0] _T_620; // @[RVC.scala 114:23:chipyard.TestHarness.RocketConfig.fir@243020.4]
  wire [25:0] _T_629; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243029.4]
  wire [28:0] _T_645; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243050.4]
  wire [27:0] _T_660; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243070.4]
  wire [28:0] _T_675; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243090.4]
  wire [24:0] _T_685; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243105.4]
  wire [24:0] _T_696; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243121.4]
  wire [24:0] _T_707; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243137.4]
  wire [24:0] _T_709; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243139.4]
  wire [24:0] _T_712; // @[RVC.scala 135:33:chipyard.TestHarness.RocketConfig.fir@243142.4]
  wire  _T_718; // @[RVC.scala 136:27:chipyard.TestHarness.RocketConfig.fir@243153.4]
  wire [31:0] _T_689_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243109.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243110.4]
  wire [31:0] _T_716_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243146.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243147.4]
  wire [31:0] _T_719_bits; // @[RVC.scala 136:22:chipyard.TestHarness.RocketConfig.fir@243154.4]
  wire [4:0] _T_719_rd; // @[RVC.scala 136:22:chipyard.TestHarness.RocketConfig.fir@243154.4]
  wire [4:0] _T_719_rs1; // @[RVC.scala 136:22:chipyard.TestHarness.RocketConfig.fir@243154.4]
  wire [4:0] _T_719_rs2; // @[RVC.scala 136:22:chipyard.TestHarness.RocketConfig.fir@243154.4]
  wire [4:0] _T_719_rs3; // @[RVC.scala 136:22:chipyard.TestHarness.RocketConfig.fir@243154.4]
  wire [24:0] _T_725; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243160.4]
  wire [24:0] _T_727; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243162.4]
  wire [24:0] _T_728; // @[RVC.scala 138:46:chipyard.TestHarness.RocketConfig.fir@243163.4]
  wire [24:0] _T_731; // @[RVC.scala 139:33:chipyard.TestHarness.RocketConfig.fir@243166.4]
  wire [31:0] _T_701_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243126.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243127.4]
  wire [31:0] _T_735_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243170.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243171.4]
  wire [31:0] _T_738_bits; // @[RVC.scala 140:25:chipyard.TestHarness.RocketConfig.fir@243178.4]
  wire [4:0] _T_738_rd; // @[RVC.scala 140:25:chipyard.TestHarness.RocketConfig.fir@243178.4]
  wire [4:0] _T_738_rs1; // @[RVC.scala 140:25:chipyard.TestHarness.RocketConfig.fir@243178.4]
  wire [31:0] _T_740_bits; // @[RVC.scala 141:10:chipyard.TestHarness.RocketConfig.fir@243180.4]
  wire [4:0] _T_740_rd; // @[RVC.scala 141:10:chipyard.TestHarness.RocketConfig.fir@243180.4]
  wire [4:0] _T_740_rs1; // @[RVC.scala 141:10:chipyard.TestHarness.RocketConfig.fir@243180.4]
  wire [4:0] _T_740_rs2; // @[RVC.scala 141:10:chipyard.TestHarness.RocketConfig.fir@243180.4]
  wire [4:0] _T_740_rs3; // @[RVC.scala 141:10:chipyard.TestHarness.RocketConfig.fir@243180.4]
  wire [8:0] _T_744; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243184.4]
  wire [28:0] _T_756; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243196.4]
  wire [7:0] _T_764; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243209.4]
  wire [27:0] _T_776; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243221.4]
  wire [28:0] _T_796; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243246.4]
  wire [4:0] _T_843; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243338.4]
  wire  _T_844; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243339.4]
  wire [31:0] _T_44_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242364.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242365.4]
  wire [31:0] _T_24_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242339.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242340.4]
  wire [31:0] _T_845_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243340.4]
  wire [4:0] _T_845_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243340.4]
  wire [4:0] _T_845_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243340.4]
  wire [4:0] _T_845_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243340.4]
  wire  _T_846; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243341.4]
  wire [31:0] _T_66_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242391.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242392.4]
  wire [31:0] _T_847_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243342.4]
  wire [4:0] _T_847_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243342.4]
  wire [4:0] _T_847_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243342.4]
  wire [4:0] _T_847_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243342.4]
  wire  _T_848; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243343.4]
  wire [31:0] _T_86_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242416.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242417.4]
  wire [31:0] _T_849_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243344.4]
  wire [4:0] _T_849_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243344.4]
  wire [4:0] _T_849_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243344.4]
  wire [4:0] _T_849_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243344.4]
  wire  _T_850; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243345.4]
  wire [31:0] _T_117_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242452.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242453.4]
  wire [31:0] _T_851_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243346.4]
  wire [4:0] _T_851_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243346.4]
  wire [4:0] _T_851_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243346.4]
  wire [4:0] _T_851_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243346.4]
  wire  _T_852; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243347.4]
  wire [31:0] _T_144_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242484.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242485.4]
  wire [31:0] _T_853_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243348.4]
  wire [4:0] _T_853_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243348.4]
  wire [4:0] _T_853_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243348.4]
  wire [4:0] _T_853_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243348.4]
  wire  _T_854; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243349.4]
  wire [31:0] _T_175_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242520.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242521.4]
  wire [31:0] _T_855_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243350.4]
  wire [4:0] _T_855_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243350.4]
  wire [4:0] _T_855_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243350.4]
  wire [4:0] _T_855_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243350.4]
  wire  _T_856; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243351.4]
  wire [31:0] _T_202_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242552.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242553.4]
  wire [31:0] _T_857_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243352.4]
  wire [4:0] _T_857_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243352.4]
  wire [4:0] _T_857_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243352.4]
  wire [4:0] _T_857_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243352.4]
  wire  _T_858; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243353.4]
  wire [31:0] _T_859_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243354.4]
  wire [4:0] _T_859_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243354.4]
  wire [4:0] _T_859_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243354.4]
  wire [4:0] _T_859_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243354.4]
  wire [4:0] _T_859_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243354.4]
  wire  _T_860; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243355.4]
  wire [31:0] _T_861_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243356.4]
  wire [4:0] _T_861_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243356.4]
  wire [4:0] _T_861_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243356.4]
  wire [4:0] _T_861_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243356.4]
  wire [4:0] _T_861_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243356.4]
  wire  _T_862; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243357.4]
  wire [31:0] _T_863_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243358.4]
  wire [4:0] _T_863_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243358.4]
  wire [4:0] _T_863_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243358.4]
  wire [4:0] _T_863_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243358.4]
  wire [4:0] _T_863_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243358.4]
  wire  _T_864; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243359.4]
  wire [31:0] _T_865_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243360.4]
  wire [4:0] _T_865_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243360.4]
  wire [4:0] _T_865_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243360.4]
  wire [4:0] _T_865_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243360.4]
  wire [4:0] _T_865_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243360.4]
  wire  _T_866; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243361.4]
  wire [31:0] _T_867_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243362.4]
  wire [4:0] _T_867_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243362.4]
  wire [4:0] _T_867_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243362.4]
  wire [4:0] _T_867_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243362.4]
  wire [4:0] _T_867_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243362.4]
  wire  _T_868; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243363.4]
  wire [31:0] _T_869_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243364.4]
  wire [4:0] _T_869_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243364.4]
  wire [4:0] _T_869_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243364.4]
  wire [4:0] _T_869_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243364.4]
  wire [4:0] _T_869_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243364.4]
  wire  _T_870; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243365.4]
  wire [31:0] _T_871_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243366.4]
  wire [4:0] _T_871_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243366.4]
  wire [4:0] _T_871_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243366.4]
  wire [4:0] _T_871_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243366.4]
  wire [4:0] _T_871_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243366.4]
  wire  _T_872; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243367.4]
  wire [31:0] _T_873_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243368.4]
  wire [4:0] _T_873_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243368.4]
  wire [4:0] _T_873_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243368.4]
  wire [4:0] _T_873_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243368.4]
  wire [4:0] _T_873_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243368.4]
  wire  _T_874; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243369.4]
  wire [31:0] _T_634_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243034.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243035.4]
  wire [31:0] _T_875_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243370.4]
  wire [4:0] _T_875_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243370.4]
  wire [4:0] _T_875_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243370.4]
  wire [4:0] _T_875_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243370.4]
  wire [4:0] _T_875_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243370.4]
  wire  _T_876; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243371.4]
  wire [31:0] _T_649_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243054.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243055.4]
  wire [31:0] _T_877_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243372.4]
  wire [4:0] _T_877_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243372.4]
  wire [4:0] _T_877_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243372.4]
  wire [4:0] _T_877_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243372.4]
  wire [4:0] _T_877_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243372.4]
  wire  _T_878; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243373.4]
  wire [31:0] _T_664_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243074.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243075.4]
  wire [31:0] _T_879_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243374.4]
  wire [4:0] _T_879_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243374.4]
  wire [4:0] _T_879_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243374.4]
  wire [4:0] _T_879_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243374.4]
  wire [4:0] _T_879_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243374.4]
  wire  _T_880; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243375.4]
  wire [31:0] _T_679_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243094.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243095.4]
  wire [31:0] _T_881_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243376.4]
  wire [4:0] _T_881_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243376.4]
  wire [4:0] _T_881_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243376.4]
  wire [4:0] _T_881_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243376.4]
  wire [4:0] _T_881_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243376.4]
  wire  _T_882; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243377.4]
  wire [31:0] _T_883_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243378.4]
  wire [4:0] _T_883_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243378.4]
  wire [4:0] _T_883_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243378.4]
  wire [4:0] _T_883_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243378.4]
  wire [4:0] _T_883_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243378.4]
  wire  _T_884; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243379.4]
  wire [31:0] _T_760_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243200.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243201.4]
  wire [31:0] _T_885_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243380.4]
  wire [4:0] _T_885_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243380.4]
  wire [4:0] _T_885_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243380.4]
  wire [4:0] _T_885_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243380.4]
  wire [4:0] _T_885_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243380.4]
  wire  _T_886; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243381.4]
  wire [31:0] _T_780_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243225.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243226.4]
  wire [31:0] _T_887_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243382.4]
  wire [4:0] _T_887_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243382.4]
  wire [4:0] _T_887_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243382.4]
  wire [4:0] _T_887_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243382.4]
  wire [4:0] _T_887_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243382.4]
  wire  _T_888; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243383.4]
  wire [31:0] _T_800_bits; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243250.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243251.4]
  wire [31:0] _T_889_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243384.4]
  wire [4:0] _T_889_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243384.4]
  wire [4:0] _T_889_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243384.4]
  wire [4:0] _T_889_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243384.4]
  wire [4:0] _T_889_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243384.4]
  wire  _T_890; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243385.4]
  wire [31:0] _T_891_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243386.4]
  wire [4:0] _T_891_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243386.4]
  wire [4:0] _T_891_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243386.4]
  wire [4:0] _T_891_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243386.4]
  wire [4:0] _T_891_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243386.4]
  wire  _T_892; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243387.4]
  wire [31:0] _T_893_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243388.4]
  wire [4:0] _T_893_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243388.4]
  wire [4:0] _T_893_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243388.4]
  wire [4:0] _T_893_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243388.4]
  wire [4:0] _T_893_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243388.4]
  wire  _T_894; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243389.4]
  wire [31:0] _T_895_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243390.4]
  wire [4:0] _T_895_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243390.4]
  wire [4:0] _T_895_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243390.4]
  wire [4:0] _T_895_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243390.4]
  wire [4:0] _T_895_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243390.4]
  wire  _T_896; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243391.4]
  wire [31:0] _T_897_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243392.4]
  wire [4:0] _T_897_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243392.4]
  wire [4:0] _T_897_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243392.4]
  wire [4:0] _T_897_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243392.4]
  wire [4:0] _T_897_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243392.4]
  wire  _T_898; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243393.4]
  wire [31:0] _T_899_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243394.4]
  wire [4:0] _T_899_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243394.4]
  wire [4:0] _T_899_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243394.4]
  wire [4:0] _T_899_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243394.4]
  wire [4:0] _T_899_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243394.4]
  wire  _T_900; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243395.4]
  wire [31:0] _T_901_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243396.4]
  wire [4:0] _T_901_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243396.4]
  wire [4:0] _T_901_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243396.4]
  wire [4:0] _T_901_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243396.4]
  wire [4:0] _T_901_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243396.4]
  wire  _T_902; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243397.4]
  wire [31:0] _T_903_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243398.4]
  wire [4:0] _T_903_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243398.4]
  wire [4:0] _T_903_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243398.4]
  wire [4:0] _T_903_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243398.4]
  wire [4:0] _T_903_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243398.4]
  wire  _T_904; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243399.4]
  assign _T_3 = |io_in[12:5]; // @[RVC.scala 54:29:chipyard.TestHarness.RocketConfig.fir@242318.4]
  assign _T_4 = _T_3 ? 7'h13 : 7'h1f; // @[RVC.scala 54:20:chipyard.TestHarness.RocketConfig.fir@242319.4]
  assign _T_14 = {2'h1,io_in[4:2]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242329.4]
  assign _T_18 = {io_in[10:7],io_in[12:11],io_in[5],io_in[6],2'h0,5'h2,3'h0,2'h1,io_in[4:2],_T_4}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242333.4]
  assign _T_28 = {io_in[6:5],io_in[12:10],3'h0}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242348.4]
  assign _T_30 = {2'h1,io_in[9:7]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242350.4]
  assign _T_36 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h7}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242356.4]
  assign _T_50 = {io_in[5],io_in[12:10],io_in[6],2'h0}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242375.4]
  assign _T_58 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h3}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242383.4]
  assign _T_78 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h3}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242408.4]
  assign _T_109 = {_T_50[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_T_50[4:0],7'h3f}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242444.4]
  assign _T_136 = {_T_28[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_T_28[4:0],7'h27}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242476.4]
  assign _T_167 = {_T_50[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_T_50[4:0],7'h23}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242512.4]
  assign _T_194 = {_T_28[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_T_28[4:0],7'h23}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242544.4]
  assign _T_205 = io_in[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@242560.4]
  assign _T_207 = {_T_205,io_in[6:2]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242562.4]
  assign _T_213 = {_T_205,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h13}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242568.4]
  assign _T_221 = |io_in[11:7]; // @[RVC.scala 78:24:chipyard.TestHarness.RocketConfig.fir@242581.4]
  assign _T_222 = _T_221 ? 7'h1b : 7'h1f; // @[RVC.scala 78:20:chipyard.TestHarness.RocketConfig.fir@242582.4]
  assign _T_233 = {_T_205,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],_T_222}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242593.4]
  assign _T_249 = {_T_205,io_in[6:2],5'h0,3'h0,io_in[11:7],7'h13}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242614.4]
  assign _T_260 = |_T_207; // @[RVC.scala 91:29:chipyard.TestHarness.RocketConfig.fir@242630.4]
  assign _T_261 = _T_260 ? 7'h37 : 7'h3f; // @[RVC.scala 91:20:chipyard.TestHarness.RocketConfig.fir@242631.4]
  assign _T_264 = io_in[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@242634.4]
  assign _T_267 = {_T_264,io_in[6:2],12'h0}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242637.4]
  assign _T_271 = {_T_267[31:12],io_in[11:7],_T_261}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242641.4]
  assign _T_279 = io_in[11:7] == 5'h0; // @[RVC.scala 93:14:chipyard.TestHarness.RocketConfig.fir@242654.4]
  assign _T_281 = io_in[11:7] == 5'h2; // @[RVC.scala 93:27:chipyard.TestHarness.RocketConfig.fir@242656.4]
  assign _T_282 = _T_279 | _T_281; // @[RVC.scala 93:21:chipyard.TestHarness.RocketConfig.fir@242657.4]
  assign _T_289 = _T_260 ? 7'h13 : 7'h1f; // @[RVC.scala 87:20:chipyard.TestHarness.RocketConfig.fir@242664.4]
  assign _T_292 = io_in[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@242667.4]
  assign _T_307 = {_T_292,io_in[4:3],io_in[5],io_in[2],io_in[6],4'h0,io_in[11:7],3'h0,io_in[11:7],_T_289}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242682.4]
  assign _T_314_bits = _T_282 ? _T_307 : _T_271; // @[RVC.scala 93:10:chipyard.TestHarness.RocketConfig.fir@242694.4]
  assign _T_314_rd = _T_282 ? io_in[11:7] : io_in[11:7]; // @[RVC.scala 93:10:chipyard.TestHarness.RocketConfig.fir@242694.4]
  assign _T_314_rs2 = _T_282 ? _T_14 : _T_14; // @[RVC.scala 93:10:chipyard.TestHarness.RocketConfig.fir@242694.4]
  assign _T_314_rs3 = _T_282 ? io_in[31:27] : io_in[31:27]; // @[RVC.scala 93:10:chipyard.TestHarness.RocketConfig.fir@242694.4]
  assign _T_325 = {io_in[12],io_in[6:2],2'h1,io_in[9:7],3'h5,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242705.4]
  assign _GEN_0 = {{5'd0}, _T_325}; // @[RVC.scala 100:23:chipyard.TestHarness.RocketConfig.fir@242717.4]
  assign _T_337 = _GEN_0 | 31'h40000000; // @[RVC.scala 100:23:chipyard.TestHarness.RocketConfig.fir@242717.4]
  assign _T_350 = {_T_205,io_in[6:2],2'h1,io_in[9:7],3'h7,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242730.4]
  assign _T_353 = {io_in[12],io_in[6:5]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242733.4]
  assign _T_354 = _T_353 == 3'h1; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242734.4]
  assign _T_355 = _T_354 ? 3'h4 : 3'h0; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242735.4]
  assign _T_356 = _T_353 == 3'h2; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242736.4]
  assign _T_357 = _T_356 ? 3'h6 : _T_355; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242737.4]
  assign _T_358 = _T_353 == 3'h3; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242738.4]
  assign _T_359 = _T_358 ? 3'h7 : _T_357; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242739.4]
  assign _T_360 = _T_353 == 3'h4; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242740.4]
  assign _T_361 = _T_360 ? 3'h0 : _T_359; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242741.4]
  assign _T_362 = _T_353 == 3'h5; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242742.4]
  assign _T_363 = _T_362 ? 3'h0 : _T_361; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242743.4]
  assign _T_364 = _T_353 == 3'h6; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242744.4]
  assign _T_365 = _T_364 ? 3'h2 : _T_363; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242745.4]
  assign _T_366 = _T_353 == 3'h7; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242746.4]
  assign _T_367 = _T_366 ? 3'h3 : _T_365; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242747.4]
  assign _T_369 = io_in[6:5] == 2'h0; // @[RVC.scala 104:30:chipyard.TestHarness.RocketConfig.fir@242749.4]
  assign _T_370 = _T_369 ? 31'h40000000 : 31'h0; // @[RVC.scala 104:22:chipyard.TestHarness.RocketConfig.fir@242750.4]
  assign _T_372 = io_in[12] ? 7'h3b : 7'h33; // @[RVC.scala 105:22:chipyard.TestHarness.RocketConfig.fir@242752.4]
  assign _T_382 = {2'h1,io_in[4:2],2'h1,io_in[9:7],_T_367,2'h1,io_in[9:7],_T_372}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242762.4]
  assign _GEN_1 = {{6'd0}, _T_382}; // @[RVC.scala 106:43:chipyard.TestHarness.RocketConfig.fir@242763.4]
  assign _T_383 = _GEN_1 | _T_370; // @[RVC.scala 106:43:chipyard.TestHarness.RocketConfig.fir@242763.4]
  assign _T_385 = io_in[11:10] == 2'h1; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242765.4]
  assign _T_386 = _T_385 ? _T_337 : {{5'd0}, _T_325}; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242766.4]
  assign _T_387 = io_in[11:10] == 2'h2; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242767.4]
  assign _T_388 = _T_387 ? _T_350 : {{1'd0}, _T_386}; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242768.4]
  assign _T_389 = io_in[11:10] == 2'h3; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@242769.4]
  assign _T_390 = _T_389 ? {{1'd0}, _T_383} : _T_388; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@242770.4]
  assign _T_401 = io_in[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@242786.4]
  assign _T_416 = {_T_401,io_in[8],io_in[10:9],io_in[6],io_in[7],io_in[2],io_in[11],io_in[5:3],1'h0}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242801.4]
  assign _T_479 = {_T_416[20],_T_416[10:1],_T_416[11],_T_416[19:12],5'h0,7'h6f}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242864.4]
  assign _T_488 = io_in[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@242878.4]
  assign _T_497 = {_T_488,io_in[6:5],io_in[2],io_in[11:10],io_in[4:3],1'h0}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242887.4]
  assign _T_546 = {_T_497[12],_T_497[10:5],5'h0,2'h1,io_in[9:7],3'h0,_T_497[4:1],_T_497[11],7'h63}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@242936.4]
  assign _T_613 = {_T_497[12],_T_497[10:5],5'h0,2'h1,io_in[9:7],3'h1,_T_497[4:1],_T_497[11],7'h63}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243008.4]
  assign _T_620 = _T_221 ? 7'h3 : 7'h1f; // @[RVC.scala 114:23:chipyard.TestHarness.RocketConfig.fir@243020.4]
  assign _T_629 = {io_in[12],io_in[6:2],io_in[11:7],3'h1,io_in[11:7],7'h13}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243029.4]
  assign _T_645 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],7'h7}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243050.4]
  assign _T_660 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],_T_620}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243070.4]
  assign _T_675 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],_T_620}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243090.4]
  assign _T_685 = {io_in[6:2],5'h0,3'h0,io_in[11:7],7'h33}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243105.4]
  assign _T_696 = {io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h33}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243121.4]
  assign _T_707 = {io_in[6:2],io_in[11:7],3'h0,12'h67}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243137.4]
  assign _T_709 = {_T_707[24:7],7'h1f}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243139.4]
  assign _T_712 = _T_221 ? _T_707 : _T_709; // @[RVC.scala 135:33:chipyard.TestHarness.RocketConfig.fir@243142.4]
  assign _T_718 = |io_in[6:2]; // @[RVC.scala 136:27:chipyard.TestHarness.RocketConfig.fir@243153.4]
  assign _T_689_bits = {{7'd0}, _T_685}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243109.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243110.4]
  assign _T_716_bits = {{7'd0}, _T_712}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243146.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243147.4]
  assign _T_719_bits = _T_718 ? _T_689_bits : _T_716_bits; // @[RVC.scala 136:22:chipyard.TestHarness.RocketConfig.fir@243154.4]
  assign _T_719_rd = _T_718 ? io_in[11:7] : 5'h0; // @[RVC.scala 136:22:chipyard.TestHarness.RocketConfig.fir@243154.4]
  assign _T_719_rs1 = _T_718 ? 5'h0 : io_in[11:7]; // @[RVC.scala 136:22:chipyard.TestHarness.RocketConfig.fir@243154.4]
  assign _T_719_rs2 = _T_718 ? io_in[6:2] : io_in[6:2]; // @[RVC.scala 136:22:chipyard.TestHarness.RocketConfig.fir@243154.4]
  assign _T_719_rs3 = _T_718 ? io_in[31:27] : io_in[31:27]; // @[RVC.scala 136:22:chipyard.TestHarness.RocketConfig.fir@243154.4]
  assign _T_725 = {io_in[6:2],io_in[11:7],3'h0,12'he7}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243160.4]
  assign _T_727 = {_T_707[24:7],7'h73}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243162.4]
  assign _T_728 = _T_727 | 25'h100000; // @[RVC.scala 138:46:chipyard.TestHarness.RocketConfig.fir@243163.4]
  assign _T_731 = _T_221 ? _T_725 : _T_728; // @[RVC.scala 139:33:chipyard.TestHarness.RocketConfig.fir@243166.4]
  assign _T_701_bits = {{7'd0}, _T_696}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243126.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243127.4]
  assign _T_735_bits = {{7'd0}, _T_731}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243170.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243171.4]
  assign _T_738_bits = _T_718 ? _T_701_bits : _T_735_bits; // @[RVC.scala 140:25:chipyard.TestHarness.RocketConfig.fir@243178.4]
  assign _T_738_rd = _T_718 ? io_in[11:7] : 5'h1; // @[RVC.scala 140:25:chipyard.TestHarness.RocketConfig.fir@243178.4]
  assign _T_738_rs1 = _T_718 ? io_in[11:7] : io_in[11:7]; // @[RVC.scala 140:25:chipyard.TestHarness.RocketConfig.fir@243178.4]
  assign _T_740_bits = io_in[12] ? _T_738_bits : _T_719_bits; // @[RVC.scala 141:10:chipyard.TestHarness.RocketConfig.fir@243180.4]
  assign _T_740_rd = io_in[12] ? _T_738_rd : _T_719_rd; // @[RVC.scala 141:10:chipyard.TestHarness.RocketConfig.fir@243180.4]
  assign _T_740_rs1 = io_in[12] ? _T_738_rs1 : _T_719_rs1; // @[RVC.scala 141:10:chipyard.TestHarness.RocketConfig.fir@243180.4]
  assign _T_740_rs2 = io_in[12] ? _T_719_rs2 : _T_719_rs2; // @[RVC.scala 141:10:chipyard.TestHarness.RocketConfig.fir@243180.4]
  assign _T_740_rs3 = io_in[12] ? _T_719_rs3 : _T_719_rs3; // @[RVC.scala 141:10:chipyard.TestHarness.RocketConfig.fir@243180.4]
  assign _T_744 = {io_in[9:7],io_in[12:10],3'h0}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243184.4]
  assign _T_756 = {_T_744[8:5],io_in[6:2],5'h2,3'h3,_T_744[4:0],7'h27}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243196.4]
  assign _T_764 = {io_in[8:7],io_in[12:9],2'h0}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243209.4]
  assign _T_776 = {_T_764[7:5],io_in[6:2],5'h2,3'h2,_T_764[4:0],7'h23}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243221.4]
  assign _T_796 = {_T_744[8:5],io_in[6:2],5'h2,3'h3,_T_744[4:0],7'h23}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243246.4]
  assign _T_843 = {io_in[1:0],io_in[15:13]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@243338.4]
  assign _T_844 = _T_843 == 5'h1; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243339.4]
  assign _T_44_bits = {{4'd0}, _T_36}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242364.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242365.4]
  assign _T_24_bits = {{2'd0}, _T_18}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242339.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242340.4]
  assign _T_845_bits = _T_844 ? _T_44_bits : _T_24_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243340.4]
  assign _T_845_rd = _T_844 ? _T_14 : _T_14; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243340.4]
  assign _T_845_rs1 = _T_844 ? _T_30 : 5'h2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243340.4]
  assign _T_845_rs3 = _T_844 ? io_in[31:27] : io_in[31:27]; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243340.4]
  assign _T_846 = _T_843 == 5'h2; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243341.4]
  assign _T_66_bits = {{5'd0}, _T_58}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242391.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242392.4]
  assign _T_847_bits = _T_846 ? _T_66_bits : _T_845_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243342.4]
  assign _T_847_rd = _T_846 ? _T_14 : _T_845_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243342.4]
  assign _T_847_rs1 = _T_846 ? _T_30 : _T_845_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243342.4]
  assign _T_847_rs3 = _T_846 ? io_in[31:27] : _T_845_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243342.4]
  assign _T_848 = _T_843 == 5'h3; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243343.4]
  assign _T_86_bits = {{4'd0}, _T_78}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242416.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242417.4]
  assign _T_849_bits = _T_848 ? _T_86_bits : _T_847_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243344.4]
  assign _T_849_rd = _T_848 ? _T_14 : _T_847_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243344.4]
  assign _T_849_rs1 = _T_848 ? _T_30 : _T_847_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243344.4]
  assign _T_849_rs3 = _T_848 ? io_in[31:27] : _T_847_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243344.4]
  assign _T_850 = _T_843 == 5'h4; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243345.4]
  assign _T_117_bits = {{5'd0}, _T_109}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242452.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242453.4]
  assign _T_851_bits = _T_850 ? _T_117_bits : _T_849_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243346.4]
  assign _T_851_rd = _T_850 ? _T_14 : _T_849_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243346.4]
  assign _T_851_rs1 = _T_850 ? _T_30 : _T_849_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243346.4]
  assign _T_851_rs3 = _T_850 ? io_in[31:27] : _T_849_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243346.4]
  assign _T_852 = _T_843 == 5'h5; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243347.4]
  assign _T_144_bits = {{4'd0}, _T_136}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242484.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242485.4]
  assign _T_853_bits = _T_852 ? _T_144_bits : _T_851_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243348.4]
  assign _T_853_rd = _T_852 ? _T_14 : _T_851_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243348.4]
  assign _T_853_rs1 = _T_852 ? _T_30 : _T_851_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243348.4]
  assign _T_853_rs3 = _T_852 ? io_in[31:27] : _T_851_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243348.4]
  assign _T_854 = _T_843 == 5'h6; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243349.4]
  assign _T_175_bits = {{5'd0}, _T_167}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242520.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242521.4]
  assign _T_855_bits = _T_854 ? _T_175_bits : _T_853_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243350.4]
  assign _T_855_rd = _T_854 ? _T_14 : _T_853_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243350.4]
  assign _T_855_rs1 = _T_854 ? _T_30 : _T_853_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243350.4]
  assign _T_855_rs3 = _T_854 ? io_in[31:27] : _T_853_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243350.4]
  assign _T_856 = _T_843 == 5'h7; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243351.4]
  assign _T_202_bits = {{4'd0}, _T_194}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@242552.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@242553.4]
  assign _T_857_bits = _T_856 ? _T_202_bits : _T_855_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243352.4]
  assign _T_857_rd = _T_856 ? _T_14 : _T_855_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243352.4]
  assign _T_857_rs1 = _T_856 ? _T_30 : _T_855_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243352.4]
  assign _T_857_rs3 = _T_856 ? io_in[31:27] : _T_855_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243352.4]
  assign _T_858 = _T_843 == 5'h8; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243353.4]
  assign _T_859_bits = _T_858 ? _T_213 : _T_857_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243354.4]
  assign _T_859_rd = _T_858 ? io_in[11:7] : _T_857_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243354.4]
  assign _T_859_rs1 = _T_858 ? io_in[11:7] : _T_857_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243354.4]
  assign _T_859_rs2 = _T_858 ? _T_14 : _T_857_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243354.4]
  assign _T_859_rs3 = _T_858 ? io_in[31:27] : _T_857_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243354.4]
  assign _T_860 = _T_843 == 5'h9; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243355.4]
  assign _T_861_bits = _T_860 ? _T_233 : _T_859_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243356.4]
  assign _T_861_rd = _T_860 ? io_in[11:7] : _T_859_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243356.4]
  assign _T_861_rs1 = _T_860 ? io_in[11:7] : _T_859_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243356.4]
  assign _T_861_rs2 = _T_860 ? _T_14 : _T_859_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243356.4]
  assign _T_861_rs3 = _T_860 ? io_in[31:27] : _T_859_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243356.4]
  assign _T_862 = _T_843 == 5'ha; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243357.4]
  assign _T_863_bits = _T_862 ? _T_249 : _T_861_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243358.4]
  assign _T_863_rd = _T_862 ? io_in[11:7] : _T_861_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243358.4]
  assign _T_863_rs1 = _T_862 ? 5'h0 : _T_861_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243358.4]
  assign _T_863_rs2 = _T_862 ? _T_14 : _T_861_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243358.4]
  assign _T_863_rs3 = _T_862 ? io_in[31:27] : _T_861_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243358.4]
  assign _T_864 = _T_843 == 5'hb; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243359.4]
  assign _T_865_bits = _T_864 ? _T_314_bits : _T_863_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243360.4]
  assign _T_865_rd = _T_864 ? _T_314_rd : _T_863_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243360.4]
  assign _T_865_rs1 = _T_864 ? _T_314_rd : _T_863_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243360.4]
  assign _T_865_rs2 = _T_864 ? _T_314_rs2 : _T_863_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243360.4]
  assign _T_865_rs3 = _T_864 ? _T_314_rs3 : _T_863_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243360.4]
  assign _T_866 = _T_843 == 5'hc; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243361.4]
  assign _T_867_bits = _T_866 ? _T_390 : _T_865_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243362.4]
  assign _T_867_rd = _T_866 ? _T_30 : _T_865_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243362.4]
  assign _T_867_rs1 = _T_866 ? _T_30 : _T_865_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243362.4]
  assign _T_867_rs2 = _T_866 ? _T_14 : _T_865_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243362.4]
  assign _T_867_rs3 = _T_866 ? io_in[31:27] : _T_865_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243362.4]
  assign _T_868 = _T_843 == 5'hd; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243363.4]
  assign _T_869_bits = _T_868 ? _T_479 : _T_867_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243364.4]
  assign _T_869_rd = _T_868 ? 5'h0 : _T_867_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243364.4]
  assign _T_869_rs1 = _T_868 ? _T_30 : _T_867_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243364.4]
  assign _T_869_rs2 = _T_868 ? _T_14 : _T_867_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243364.4]
  assign _T_869_rs3 = _T_868 ? io_in[31:27] : _T_867_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243364.4]
  assign _T_870 = _T_843 == 5'he; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243365.4]
  assign _T_871_bits = _T_870 ? _T_546 : _T_869_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243366.4]
  assign _T_871_rd = _T_870 ? _T_30 : _T_869_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243366.4]
  assign _T_871_rs1 = _T_870 ? _T_30 : _T_869_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243366.4]
  assign _T_871_rs2 = _T_870 ? 5'h0 : _T_869_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243366.4]
  assign _T_871_rs3 = _T_870 ? io_in[31:27] : _T_869_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243366.4]
  assign _T_872 = _T_843 == 5'hf; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243367.4]
  assign _T_873_bits = _T_872 ? _T_613 : _T_871_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243368.4]
  assign _T_873_rd = _T_872 ? 5'h0 : _T_871_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243368.4]
  assign _T_873_rs1 = _T_872 ? _T_30 : _T_871_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243368.4]
  assign _T_873_rs2 = _T_872 ? 5'h0 : _T_871_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243368.4]
  assign _T_873_rs3 = _T_872 ? io_in[31:27] : _T_871_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243368.4]
  assign _T_874 = _T_843 == 5'h10; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243369.4]
  assign _T_634_bits = {{6'd0}, _T_629}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243034.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243035.4]
  assign _T_875_bits = _T_874 ? _T_634_bits : _T_873_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243370.4]
  assign _T_875_rd = _T_874 ? io_in[11:7] : _T_873_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243370.4]
  assign _T_875_rs1 = _T_874 ? io_in[11:7] : _T_873_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243370.4]
  assign _T_875_rs2 = _T_874 ? io_in[6:2] : _T_873_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243370.4]
  assign _T_875_rs3 = _T_874 ? io_in[31:27] : _T_873_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243370.4]
  assign _T_876 = _T_843 == 5'h11; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243371.4]
  assign _T_649_bits = {{3'd0}, _T_645}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243054.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243055.4]
  assign _T_877_bits = _T_876 ? _T_649_bits : _T_875_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243372.4]
  assign _T_877_rd = _T_876 ? io_in[11:7] : _T_875_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243372.4]
  assign _T_877_rs1 = _T_876 ? 5'h2 : _T_875_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243372.4]
  assign _T_877_rs2 = _T_876 ? io_in[6:2] : _T_875_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243372.4]
  assign _T_877_rs3 = _T_876 ? io_in[31:27] : _T_875_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243372.4]
  assign _T_878 = _T_843 == 5'h12; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243373.4]
  assign _T_664_bits = {{4'd0}, _T_660}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243074.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243075.4]
  assign _T_879_bits = _T_878 ? _T_664_bits : _T_877_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243374.4]
  assign _T_879_rd = _T_878 ? io_in[11:7] : _T_877_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243374.4]
  assign _T_879_rs1 = _T_878 ? 5'h2 : _T_877_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243374.4]
  assign _T_879_rs2 = _T_878 ? io_in[6:2] : _T_877_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243374.4]
  assign _T_879_rs3 = _T_878 ? io_in[31:27] : _T_877_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243374.4]
  assign _T_880 = _T_843 == 5'h13; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243375.4]
  assign _T_679_bits = {{3'd0}, _T_675}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243094.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243095.4]
  assign _T_881_bits = _T_880 ? _T_679_bits : _T_879_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243376.4]
  assign _T_881_rd = _T_880 ? io_in[11:7] : _T_879_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243376.4]
  assign _T_881_rs1 = _T_880 ? 5'h2 : _T_879_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243376.4]
  assign _T_881_rs2 = _T_880 ? io_in[6:2] : _T_879_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243376.4]
  assign _T_881_rs3 = _T_880 ? io_in[31:27] : _T_879_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243376.4]
  assign _T_882 = _T_843 == 5'h14; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243377.4]
  assign _T_883_bits = _T_882 ? _T_740_bits : _T_881_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243378.4]
  assign _T_883_rd = _T_882 ? _T_740_rd : _T_881_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243378.4]
  assign _T_883_rs1 = _T_882 ? _T_740_rs1 : _T_881_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243378.4]
  assign _T_883_rs2 = _T_882 ? _T_740_rs2 : _T_881_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243378.4]
  assign _T_883_rs3 = _T_882 ? _T_740_rs3 : _T_881_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243378.4]
  assign _T_884 = _T_843 == 5'h15; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243379.4]
  assign _T_760_bits = {{3'd0}, _T_756}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243200.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243201.4]
  assign _T_885_bits = _T_884 ? _T_760_bits : _T_883_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243380.4]
  assign _T_885_rd = _T_884 ? io_in[11:7] : _T_883_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243380.4]
  assign _T_885_rs1 = _T_884 ? 5'h2 : _T_883_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243380.4]
  assign _T_885_rs2 = _T_884 ? io_in[6:2] : _T_883_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243380.4]
  assign _T_885_rs3 = _T_884 ? io_in[31:27] : _T_883_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243380.4]
  assign _T_886 = _T_843 == 5'h16; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243381.4]
  assign _T_780_bits = {{4'd0}, _T_776}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243225.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243226.4]
  assign _T_887_bits = _T_886 ? _T_780_bits : _T_885_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243382.4]
  assign _T_887_rd = _T_886 ? io_in[11:7] : _T_885_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243382.4]
  assign _T_887_rs1 = _T_886 ? 5'h2 : _T_885_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243382.4]
  assign _T_887_rs2 = _T_886 ? io_in[6:2] : _T_885_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243382.4]
  assign _T_887_rs3 = _T_886 ? io_in[31:27] : _T_885_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243382.4]
  assign _T_888 = _T_843 == 5'h17; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243383.4]
  assign _T_800_bits = {{3'd0}, _T_796}; // @[RVC.scala 22:19:chipyard.TestHarness.RocketConfig.fir@243250.4 RVC.scala 23:14:chipyard.TestHarness.RocketConfig.fir@243251.4]
  assign _T_889_bits = _T_888 ? _T_800_bits : _T_887_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243384.4]
  assign _T_889_rd = _T_888 ? io_in[11:7] : _T_887_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243384.4]
  assign _T_889_rs1 = _T_888 ? 5'h2 : _T_887_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243384.4]
  assign _T_889_rs2 = _T_888 ? io_in[6:2] : _T_887_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243384.4]
  assign _T_889_rs3 = _T_888 ? io_in[31:27] : _T_887_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243384.4]
  assign _T_890 = _T_843 == 5'h18; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243385.4]
  assign _T_891_bits = _T_890 ? io_in : _T_889_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243386.4]
  assign _T_891_rd = _T_890 ? io_in[11:7] : _T_889_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243386.4]
  assign _T_891_rs1 = _T_890 ? io_in[19:15] : _T_889_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243386.4]
  assign _T_891_rs2 = _T_890 ? io_in[24:20] : _T_889_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243386.4]
  assign _T_891_rs3 = _T_890 ? io_in[31:27] : _T_889_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243386.4]
  assign _T_892 = _T_843 == 5'h19; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243387.4]
  assign _T_893_bits = _T_892 ? io_in : _T_891_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243388.4]
  assign _T_893_rd = _T_892 ? io_in[11:7] : _T_891_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243388.4]
  assign _T_893_rs1 = _T_892 ? io_in[19:15] : _T_891_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243388.4]
  assign _T_893_rs2 = _T_892 ? io_in[24:20] : _T_891_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243388.4]
  assign _T_893_rs3 = _T_892 ? io_in[31:27] : _T_891_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243388.4]
  assign _T_894 = _T_843 == 5'h1a; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243389.4]
  assign _T_895_bits = _T_894 ? io_in : _T_893_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243390.4]
  assign _T_895_rd = _T_894 ? io_in[11:7] : _T_893_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243390.4]
  assign _T_895_rs1 = _T_894 ? io_in[19:15] : _T_893_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243390.4]
  assign _T_895_rs2 = _T_894 ? io_in[24:20] : _T_893_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243390.4]
  assign _T_895_rs3 = _T_894 ? io_in[31:27] : _T_893_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243390.4]
  assign _T_896 = _T_843 == 5'h1b; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243391.4]
  assign _T_897_bits = _T_896 ? io_in : _T_895_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243392.4]
  assign _T_897_rd = _T_896 ? io_in[11:7] : _T_895_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243392.4]
  assign _T_897_rs1 = _T_896 ? io_in[19:15] : _T_895_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243392.4]
  assign _T_897_rs2 = _T_896 ? io_in[24:20] : _T_895_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243392.4]
  assign _T_897_rs3 = _T_896 ? io_in[31:27] : _T_895_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243392.4]
  assign _T_898 = _T_843 == 5'h1c; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243393.4]
  assign _T_899_bits = _T_898 ? io_in : _T_897_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243394.4]
  assign _T_899_rd = _T_898 ? io_in[11:7] : _T_897_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243394.4]
  assign _T_899_rs1 = _T_898 ? io_in[19:15] : _T_897_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243394.4]
  assign _T_899_rs2 = _T_898 ? io_in[24:20] : _T_897_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243394.4]
  assign _T_899_rs3 = _T_898 ? io_in[31:27] : _T_897_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243394.4]
  assign _T_900 = _T_843 == 5'h1d; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243395.4]
  assign _T_901_bits = _T_900 ? io_in : _T_899_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243396.4]
  assign _T_901_rd = _T_900 ? io_in[11:7] : _T_899_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243396.4]
  assign _T_901_rs1 = _T_900 ? io_in[19:15] : _T_899_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243396.4]
  assign _T_901_rs2 = _T_900 ? io_in[24:20] : _T_899_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243396.4]
  assign _T_901_rs3 = _T_900 ? io_in[31:27] : _T_899_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243396.4]
  assign _T_902 = _T_843 == 5'h1e; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243397.4]
  assign _T_903_bits = _T_902 ? io_in : _T_901_bits; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243398.4]
  assign _T_903_rd = _T_902 ? io_in[11:7] : _T_901_rd; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243398.4]
  assign _T_903_rs1 = _T_902 ? io_in[19:15] : _T_901_rs1; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243398.4]
  assign _T_903_rs2 = _T_902 ? io_in[24:20] : _T_901_rs2; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243398.4]
  assign _T_903_rs3 = _T_902 ? io_in[31:27] : _T_901_rs3; // @[package.scala 32:76:chipyard.TestHarness.RocketConfig.fir@243398.4]
  assign _T_904 = _T_843 == 5'h1f; // @[package.scala 32:86:chipyard.TestHarness.RocketConfig.fir@243399.4]
  assign io_out_bits = _T_904 ? io_in : _T_903_bits; // @[RVC.scala 165:12:chipyard.TestHarness.RocketConfig.fir@243405.4]
  assign io_out_rd = _T_904 ? io_in[11:7] : _T_903_rd; // @[RVC.scala 165:12:chipyard.TestHarness.RocketConfig.fir@243404.4]
  assign io_out_rs1 = _T_904 ? io_in[19:15] : _T_903_rs1; // @[RVC.scala 165:12:chipyard.TestHarness.RocketConfig.fir@243403.4]
  assign io_out_rs2 = _T_904 ? io_in[24:20] : _T_903_rs2; // @[RVC.scala 165:12:chipyard.TestHarness.RocketConfig.fir@243402.4]
  assign io_out_rs3 = _T_904 ? io_in[31:27] : _T_903_rs3; // @[RVC.scala 165:12:chipyard.TestHarness.RocketConfig.fir@243401.4]
  assign io_rvc = io_in[1:0] != 2'h3; // @[RVC.scala 164:12:chipyard.TestHarness.RocketConfig.fir@242316.4]
endmodule
