module package_Anon_117( // @[:chipyard.TestHarness.RocketConfig.fir@240846.2]
  input  [2:0] io_x, // @[:chipyard.TestHarness.RocketConfig.fir@240849.4]
  output [2:0] io_y // @[:chipyard.TestHarness.RocketConfig.fir@240849.4]
);
  assign io_y = io_x; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@240854.4]
endmodule
