module TLB_1( // @[:chipyard.TestHarness.RocketConfig.fir@220830.2]
  input         clock, // @[:chipyard.TestHarness.RocketConfig.fir@220831.4]
  input         reset, // @[:chipyard.TestHarness.RocketConfig.fir@220832.4]
  output        io_req_ready, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_req_valid, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [39:0] io_req_bits_vaddr, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  output        io_resp_miss, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  output [31:0] io_resp_paddr, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  output        io_resp_pf_inst, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  output        io_resp_ae_inst, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  output        io_resp_cacheable, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_sfence_valid, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_sfence_bits_rs1, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_sfence_bits_rs2, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [38:0] io_sfence_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_req_ready, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  output        io_ptw_req_valid, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  output        io_ptw_req_bits_valid, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  output [26:0] io_ptw_req_bits_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_resp_valid, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_resp_bits_ae, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [53:0] io_ptw_resp_bits_pte_ppn, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_resp_bits_pte_d, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_resp_bits_pte_a, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_resp_bits_pte_g, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_resp_bits_pte_u, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_resp_bits_pte_x, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_resp_bits_pte_w, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_resp_bits_pte_r, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_resp_bits_pte_v, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [1:0]  io_ptw_resp_bits_level, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_resp_bits_homogeneous, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [3:0]  io_ptw_ptbr_mode, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_status_debug, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [1:0]  io_ptw_status_prv, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_0_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [1:0]  io_ptw_pmp_0_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_0_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_0_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_0_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [29:0] io_ptw_pmp_0_addr, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [31:0] io_ptw_pmp_0_mask, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_1_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [1:0]  io_ptw_pmp_1_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_1_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_1_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_1_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [29:0] io_ptw_pmp_1_addr, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [31:0] io_ptw_pmp_1_mask, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_2_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [1:0]  io_ptw_pmp_2_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_2_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_2_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_2_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [29:0] io_ptw_pmp_2_addr, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [31:0] io_ptw_pmp_2_mask, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_3_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [1:0]  io_ptw_pmp_3_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_3_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_3_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_3_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [29:0] io_ptw_pmp_3_addr, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [31:0] io_ptw_pmp_3_mask, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_4_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [1:0]  io_ptw_pmp_4_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_4_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_4_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_4_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [29:0] io_ptw_pmp_4_addr, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [31:0] io_ptw_pmp_4_mask, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_5_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [1:0]  io_ptw_pmp_5_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_5_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_5_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_5_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [29:0] io_ptw_pmp_5_addr, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [31:0] io_ptw_pmp_5_mask, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_6_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [1:0]  io_ptw_pmp_6_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_6_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_6_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_6_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [29:0] io_ptw_pmp_6_addr, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [31:0] io_ptw_pmp_6_mask, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_7_cfg_l, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [1:0]  io_ptw_pmp_7_cfg_a, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_7_cfg_x, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_7_cfg_w, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_ptw_pmp_7_cfg_r, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [29:0] io_ptw_pmp_7_addr, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input  [31:0] io_ptw_pmp_7_mask, // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
  input         io_kill // @[:chipyard.TestHarness.RocketConfig.fir@220833.4]
);
  wire [19:0] package_Anon_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire [19:0] package_Anon_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire  package_Anon_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
  wire [1:0] pmp_io_prv; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_0_cfg_l; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_0_cfg_x; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_0_cfg_w; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_0_cfg_r; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [29:0] pmp_io_pmp_0_addr; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [31:0] pmp_io_pmp_0_mask; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_1_cfg_l; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_1_cfg_x; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_1_cfg_w; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_1_cfg_r; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [29:0] pmp_io_pmp_1_addr; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [31:0] pmp_io_pmp_1_mask; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_2_cfg_l; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_2_cfg_x; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_2_cfg_w; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_2_cfg_r; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [29:0] pmp_io_pmp_2_addr; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [31:0] pmp_io_pmp_2_mask; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_3_cfg_l; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_3_cfg_x; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_3_cfg_w; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_3_cfg_r; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [29:0] pmp_io_pmp_3_addr; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [31:0] pmp_io_pmp_3_mask; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_4_cfg_l; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_4_cfg_x; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_4_cfg_w; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_4_cfg_r; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [29:0] pmp_io_pmp_4_addr; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [31:0] pmp_io_pmp_4_mask; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_5_cfg_l; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_5_cfg_x; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_5_cfg_w; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_5_cfg_r; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [29:0] pmp_io_pmp_5_addr; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [31:0] pmp_io_pmp_5_mask; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_6_cfg_l; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_6_cfg_x; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_6_cfg_w; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_6_cfg_r; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [29:0] pmp_io_pmp_6_addr; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [31:0] pmp_io_pmp_6_mask; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_7_cfg_l; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_7_cfg_x; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_7_cfg_w; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_pmp_7_cfg_r; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [29:0] pmp_io_pmp_7_addr; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [31:0] pmp_io_pmp_7_mask; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [31:0] pmp_io_addr; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_r; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_w; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire  pmp_io_x; // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
  wire [19:0] package_Anon_1_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire [19:0] package_Anon_1_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire  package_Anon_1_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
  wire [19:0] package_Anon_2_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire [19:0] package_Anon_2_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire  package_Anon_2_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
  wire [19:0] package_Anon_3_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire [19:0] package_Anon_3_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire  package_Anon_3_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
  wire [19:0] package_Anon_4_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire [19:0] package_Anon_4_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire  package_Anon_4_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
  wire [19:0] package_Anon_5_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire [19:0] package_Anon_5_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire  package_Anon_5_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
  wire [19:0] package_Anon_6_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire [19:0] package_Anon_6_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire  package_Anon_6_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
  wire [19:0] package_Anon_7_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire [19:0] package_Anon_7_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire  package_Anon_7_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
  wire [19:0] package_Anon_8_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire [19:0] package_Anon_8_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire  package_Anon_8_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
  wire [19:0] package_Anon_9_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire [19:0] package_Anon_9_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire  package_Anon_9_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
  wire [19:0] package_Anon_10_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire [19:0] package_Anon_10_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire  package_Anon_10_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
  wire [19:0] package_Anon_11_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire [19:0] package_Anon_11_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire  package_Anon_11_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
  wire [19:0] package_Anon_12_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire [19:0] package_Anon_12_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire  package_Anon_12_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
  wire [19:0] package_Anon_13_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire [19:0] package_Anon_13_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire  package_Anon_13_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
  wire [19:0] package_Anon_14_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire [19:0] package_Anon_14_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire  package_Anon_14_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
  wire [19:0] package_Anon_15_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire [19:0] package_Anon_15_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire  package_Anon_15_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
  wire [19:0] package_Anon_16_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire [19:0] package_Anon_16_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire  package_Anon_16_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
  wire [19:0] package_Anon_17_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire [19:0] package_Anon_17_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire  package_Anon_17_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
  wire [19:0] package_Anon_18_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire [19:0] package_Anon_18_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire  package_Anon_18_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
  wire [19:0] package_Anon_19_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire [19:0] package_Anon_19_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire  package_Anon_19_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
  wire [19:0] package_Anon_20_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire [19:0] package_Anon_20_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire  package_Anon_20_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
  wire [19:0] package_Anon_21_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire [19:0] package_Anon_21_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire  package_Anon_21_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
  wire [19:0] package_Anon_22_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire [19:0] package_Anon_22_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire  package_Anon_22_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
  wire [19:0] package_Anon_23_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire [19:0] package_Anon_23_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire  package_Anon_23_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
  wire [19:0] package_Anon_24_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire [19:0] package_Anon_24_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire  package_Anon_24_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
  wire [19:0] package_Anon_25_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire [19:0] package_Anon_25_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire  package_Anon_25_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
  wire [19:0] package_Anon_26_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire [19:0] package_Anon_26_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire  package_Anon_26_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
  wire [19:0] package_Anon_27_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire [19:0] package_Anon_27_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire  package_Anon_27_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
  wire [19:0] package_Anon_28_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire [19:0] package_Anon_28_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire  package_Anon_28_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
  wire [19:0] package_Anon_29_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire [19:0] package_Anon_29_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire  package_Anon_29_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
  wire [19:0] package_Anon_30_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire [19:0] package_Anon_30_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire  package_Anon_30_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
  wire [19:0] package_Anon_31_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire [19:0] package_Anon_31_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire  package_Anon_31_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
  wire [19:0] package_Anon_32_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire [19:0] package_Anon_32_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire  package_Anon_32_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
  wire [19:0] package_Anon_33_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire [19:0] package_Anon_33_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire  package_Anon_33_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
  wire [19:0] package_Anon_34_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire [19:0] package_Anon_34_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire  package_Anon_34_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
  wire [19:0] package_Anon_35_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire [19:0] package_Anon_35_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire  package_Anon_35_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
  wire [19:0] package_Anon_36_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire [19:0] package_Anon_36_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire  package_Anon_36_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
  wire [19:0] package_Anon_37_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire [19:0] package_Anon_37_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire  package_Anon_37_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
  wire [19:0] package_Anon_38_io_x_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_x_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_x_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_x_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_x_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_x_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_x_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_x_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_x_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_x_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_x_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_x_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_x_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire [19:0] package_Anon_38_io_y_ppn; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_y_u; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_y_ae; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_y_sw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_y_sx; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_y_sr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_y_pw; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_y_px; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_y_pr; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_y_pal; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_y_paa; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_y_eff; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  wire  package_Anon_38_io_y_c; // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
  reg [26:0] sectored_entries_0_tag; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_0;
  reg [33:0] sectored_entries_0_data_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_1;
  reg [33:0] sectored_entries_0_data_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_2;
  reg [33:0] sectored_entries_0_data_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_3;
  reg [33:0] sectored_entries_0_data_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_4;
  reg  sectored_entries_0_valid_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_5;
  reg  sectored_entries_0_valid_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_6;
  reg  sectored_entries_0_valid_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_7;
  reg  sectored_entries_0_valid_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_8;
  reg [26:0] sectored_entries_1_tag; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_9;
  reg [33:0] sectored_entries_1_data_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_10;
  reg [33:0] sectored_entries_1_data_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_11;
  reg [33:0] sectored_entries_1_data_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_12;
  reg [33:0] sectored_entries_1_data_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_13;
  reg  sectored_entries_1_valid_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_14;
  reg  sectored_entries_1_valid_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_15;
  reg  sectored_entries_1_valid_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_16;
  reg  sectored_entries_1_valid_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_17;
  reg [26:0] sectored_entries_2_tag; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_18;
  reg [33:0] sectored_entries_2_data_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_19;
  reg [33:0] sectored_entries_2_data_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_20;
  reg [33:0] sectored_entries_2_data_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_21;
  reg [33:0] sectored_entries_2_data_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_22;
  reg  sectored_entries_2_valid_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_23;
  reg  sectored_entries_2_valid_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_24;
  reg  sectored_entries_2_valid_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_25;
  reg  sectored_entries_2_valid_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_26;
  reg [26:0] sectored_entries_3_tag; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_27;
  reg [33:0] sectored_entries_3_data_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_28;
  reg [33:0] sectored_entries_3_data_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_29;
  reg [33:0] sectored_entries_3_data_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_30;
  reg [33:0] sectored_entries_3_data_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_31;
  reg  sectored_entries_3_valid_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_32;
  reg  sectored_entries_3_valid_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_33;
  reg  sectored_entries_3_valid_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_34;
  reg  sectored_entries_3_valid_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_35;
  reg [26:0] sectored_entries_4_tag; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_36;
  reg [33:0] sectored_entries_4_data_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_37;
  reg [33:0] sectored_entries_4_data_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_38;
  reg [33:0] sectored_entries_4_data_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_39;
  reg [33:0] sectored_entries_4_data_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_40;
  reg  sectored_entries_4_valid_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_41;
  reg  sectored_entries_4_valid_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_42;
  reg  sectored_entries_4_valid_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_43;
  reg  sectored_entries_4_valid_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_44;
  reg [26:0] sectored_entries_5_tag; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_45;
  reg [33:0] sectored_entries_5_data_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_46;
  reg [33:0] sectored_entries_5_data_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_47;
  reg [33:0] sectored_entries_5_data_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_48;
  reg [33:0] sectored_entries_5_data_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_49;
  reg  sectored_entries_5_valid_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_50;
  reg  sectored_entries_5_valid_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_51;
  reg  sectored_entries_5_valid_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_52;
  reg  sectored_entries_5_valid_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_53;
  reg [26:0] sectored_entries_6_tag; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_54;
  reg [33:0] sectored_entries_6_data_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_55;
  reg [33:0] sectored_entries_6_data_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_56;
  reg [33:0] sectored_entries_6_data_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_57;
  reg [33:0] sectored_entries_6_data_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_58;
  reg  sectored_entries_6_valid_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_59;
  reg  sectored_entries_6_valid_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_60;
  reg  sectored_entries_6_valid_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_61;
  reg  sectored_entries_6_valid_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_62;
  reg [26:0] sectored_entries_7_tag; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_63;
  reg [33:0] sectored_entries_7_data_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_64;
  reg [33:0] sectored_entries_7_data_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_65;
  reg [33:0] sectored_entries_7_data_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_66;
  reg [33:0] sectored_entries_7_data_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [63:0] _RAND_67;
  reg  sectored_entries_7_valid_0; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_68;
  reg  sectored_entries_7_valid_1; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_69;
  reg  sectored_entries_7_valid_2; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_70;
  reg  sectored_entries_7_valid_3; // @[TLB.scala 161:29:chipyard.TestHarness.RocketConfig.fir@220838.4]
  reg [31:0] _RAND_71;
  reg [1:0] superpage_entries_0_level; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [31:0] _RAND_72;
  reg [26:0] superpage_entries_0_tag; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [31:0] _RAND_73;
  reg [33:0] superpage_entries_0_data_0; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [63:0] _RAND_74;
  reg  superpage_entries_0_valid_0; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [31:0] _RAND_75;
  reg [1:0] superpage_entries_1_level; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [31:0] _RAND_76;
  reg [26:0] superpage_entries_1_tag; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [31:0] _RAND_77;
  reg [33:0] superpage_entries_1_data_0; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [63:0] _RAND_78;
  reg  superpage_entries_1_valid_0; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [31:0] _RAND_79;
  reg [1:0] superpage_entries_2_level; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [31:0] _RAND_80;
  reg [26:0] superpage_entries_2_tag; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [31:0] _RAND_81;
  reg [33:0] superpage_entries_2_data_0; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [63:0] _RAND_82;
  reg  superpage_entries_2_valid_0; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [31:0] _RAND_83;
  reg [1:0] superpage_entries_3_level; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [31:0] _RAND_84;
  reg [26:0] superpage_entries_3_tag; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [31:0] _RAND_85;
  reg [33:0] superpage_entries_3_data_0; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [63:0] _RAND_86;
  reg  superpage_entries_3_valid_0; // @[TLB.scala 162:30:chipyard.TestHarness.RocketConfig.fir@220839.4]
  reg [31:0] _RAND_87;
  reg [1:0] special_entry_level; // @[TLB.scala 163:56:chipyard.TestHarness.RocketConfig.fir@220840.4]
  reg [31:0] _RAND_88;
  reg [26:0] special_entry_tag; // @[TLB.scala 163:56:chipyard.TestHarness.RocketConfig.fir@220840.4]
  reg [31:0] _RAND_89;
  reg [33:0] special_entry_data_0; // @[TLB.scala 163:56:chipyard.TestHarness.RocketConfig.fir@220840.4]
  reg [63:0] _RAND_90;
  reg  special_entry_valid_0; // @[TLB.scala 163:56:chipyard.TestHarness.RocketConfig.fir@220840.4]
  reg [31:0] _RAND_91;
  reg [1:0] state; // @[TLB.scala 168:18:chipyard.TestHarness.RocketConfig.fir@220841.4]
  reg [31:0] _RAND_92;
  reg [26:0] r_refill_tag; // @[TLB.scala 169:25:chipyard.TestHarness.RocketConfig.fir@220842.4]
  reg [31:0] _RAND_93;
  reg [1:0] r_superpage_repl_addr; // @[TLB.scala 170:34:chipyard.TestHarness.RocketConfig.fir@220843.4]
  reg [31:0] _RAND_94;
  reg [2:0] r_sectored_repl_addr; // @[TLB.scala 171:33:chipyard.TestHarness.RocketConfig.fir@220844.4]
  reg [31:0] _RAND_95;
  reg [2:0] r_sectored_hit_addr; // @[TLB.scala 172:32:chipyard.TestHarness.RocketConfig.fir@220845.4]
  reg [31:0] _RAND_96;
  reg  r_sectored_hit; // @[TLB.scala 173:27:chipyard.TestHarness.RocketConfig.fir@220846.4]
  reg [31:0] _RAND_97;
  wire  priv_s; // @[TLB.scala 176:20:chipyard.TestHarness.RocketConfig.fir@220847.4]
  wire  priv_uses_vm; // @[TLB.scala 177:27:chipyard.TestHarness.RocketConfig.fir@220848.4]
  wire  vm_enabled; // @[TLB.scala 178:83:chipyard.TestHarness.RocketConfig.fir@220851.4]
  wire [26:0] vpn; // @[TLB.scala 181:30:chipyard.TestHarness.RocketConfig.fir@220854.4]
  wire [19:0] refill_ppn; // @[TLB.scala 182:44:chipyard.TestHarness.RocketConfig.fir@220855.4]
  wire  _T_4; // @[package.scala 15:47:chipyard.TestHarness.RocketConfig.fir@220857.4]
  wire  _T_5; // @[package.scala 15:47:chipyard.TestHarness.RocketConfig.fir@220858.4]
  wire  invalidate_refill; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@220859.4]
  wire  _T_25; // @[TLB.scala 107:28:chipyard.TestHarness.RocketConfig.fir@220902.4]
  wire [26:0] _T_27; // @[TLB.scala 108:28:chipyard.TestHarness.RocketConfig.fir@220904.4]
  wire [26:0] _GEN_950; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@220905.4]
  wire [26:0] _T_28; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@220905.4]
  wire  _T_31; // @[TLB.scala 107:28:chipyard.TestHarness.RocketConfig.fir@220908.4]
  wire [26:0] _T_33; // @[TLB.scala 108:28:chipyard.TestHarness.RocketConfig.fir@220910.4]
  wire [26:0] _T_34; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@220911.4]
  wire [19:0] _T_36; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@220913.4]
  wire [27:0] _T_38; // @[TLB.scala 186:20:chipyard.TestHarness.RocketConfig.fir@220915.4]
  wire [27:0] mpu_ppn; // @[TLB.scala 185:20:chipyard.TestHarness.RocketConfig.fir@220916.4]
  wire [39:0] mpu_physaddr; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@220918.4]
  wire [2:0] _T_42; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@220921.4]
  wire [2:0] mpu_priv; // @[TLB.scala 188:27:chipyard.TestHarness.RocketConfig.fir@220922.4]
  wire [39:0] _T_43; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220938.4]
  wire [40:0] _T_44; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220939.4]
  wire [40:0] _T_46; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220941.4]
  wire  _T_47; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220942.4]
  wire [39:0] _T_48; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220943.4]
  wire [40:0] _T_49; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220944.4]
  wire [40:0] _T_51; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220946.4]
  wire  _T_52; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220947.4]
  wire [39:0] _T_53; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220948.4]
  wire [40:0] _T_54; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220949.4]
  wire [40:0] _T_56; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220951.4]
  wire  _T_57; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220952.4]
  wire [39:0] _T_58; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220953.4]
  wire [40:0] _T_59; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220954.4]
  wire [40:0] _T_61; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220956.4]
  wire  _T_62; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220957.4]
  wire [39:0] _T_63; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220958.4]
  wire [40:0] _T_64; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220959.4]
  wire [40:0] _T_66; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220961.4]
  wire  _T_67; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220962.4]
  wire [40:0] _T_69; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220964.4]
  wire [40:0] _T_71; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220966.4]
  wire  _T_72; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220967.4]
  wire [39:0] _T_73; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220968.4]
  wire [40:0] _T_74; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220969.4]
  wire [40:0] _T_76; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220971.4]
  wire  _T_77; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220972.4]
  wire [39:0] _T_78; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220973.4]
  wire [40:0] _T_79; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220974.4]
  wire [40:0] _T_81; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220976.4]
  wire  _T_82; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220977.4]
  wire  _T_84; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220988.4]
  wire  _T_85; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220989.4]
  wire  _T_86; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220990.4]
  wire  _T_87; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220991.4]
  wire  _T_88; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220992.4]
  wire  _T_89; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220993.4]
  wire  legal_address; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220994.4]
  wire [40:0] _T_98; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221003.4]
  wire  _T_99; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221004.4]
  wire  cacheable; // @[TLB.scala 196:19:chipyard.TestHarness.RocketConfig.fir@221010.4]
  wire [40:0] _T_163; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221071.4]
  wire  _T_164; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221072.4]
  wire  _T_171; // @[TLBPermissions.scala 82:66:chipyard.TestHarness.RocketConfig.fir@221079.4]
  wire  _T_192; // @[TLB.scala 199:39:chipyard.TestHarness.RocketConfig.fir@221100.4]
  wire  deny_access_to_debug; // @[TLB.scala 199:48:chipyard.TestHarness.RocketConfig.fir@221106.4]
  wire  _T_204; // @[TLB.scala 200:44:chipyard.TestHarness.RocketConfig.fir@221113.4]
  wire  _T_205; // @[TLB.scala 200:41:chipyard.TestHarness.RocketConfig.fir@221114.4]
  wire  prot_r; // @[TLB.scala 200:66:chipyard.TestHarness.RocketConfig.fir@221115.4]
  wire [40:0] _T_209; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221119.4]
  wire  _T_210; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221120.4]
  wire [40:0] _T_214; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221124.4]
  wire  _T_215; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221125.4]
  wire [39:0] _T_216; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@221126.4]
  wire [40:0] _T_217; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@221127.4]
  wire [40:0] _T_219; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221129.4]
  wire  _T_220; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221130.4]
  wire  _T_226; // @[Parameters.scala 528:89:chipyard.TestHarness.RocketConfig.fir@221136.4]
  wire  _T_227; // @[Parameters.scala 528:89:chipyard.TestHarness.RocketConfig.fir@221137.4]
  wire  _T_228; // @[Parameters.scala 528:89:chipyard.TestHarness.RocketConfig.fir@221138.4]
  wire  _T_238; // @[TLB.scala 196:19:chipyard.TestHarness.RocketConfig.fir@221149.4]
  wire  _T_240; // @[TLB.scala 201:45:chipyard.TestHarness.RocketConfig.fir@221151.4]
  wire  prot_w; // @[TLB.scala 201:70:chipyard.TestHarness.RocketConfig.fir@221152.4]
  wire  _T_337; // @[TLB.scala 196:19:chipyard.TestHarness.RocketConfig.fir@221254.4]
  wire  _T_339; // @[TLB.scala 204:40:chipyard.TestHarness.RocketConfig.fir@221256.4]
  wire  prot_x; // @[TLB.scala 204:65:chipyard.TestHarness.RocketConfig.fir@221257.4]
  wire [40:0] _T_360; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221278.4]
  wire  _T_361; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221279.4]
  wire [40:0] _T_365; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221283.4]
  wire  _T_366; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221284.4]
  wire [40:0] _T_375; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221293.4]
  wire  _T_376; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221294.4]
  wire  _T_377; // @[Parameters.scala 528:89:chipyard.TestHarness.RocketConfig.fir@221295.4]
  wire  _T_378; // @[Parameters.scala 528:89:chipyard.TestHarness.RocketConfig.fir@221296.4]
  wire  _T_379; // @[Parameters.scala 528:89:chipyard.TestHarness.RocketConfig.fir@221297.4]
  wire  prot_eff; // @[TLB.scala 196:19:chipyard.TestHarness.RocketConfig.fir@221303.4]
  wire  _T_384; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221304.4]
  wire  _T_385; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221305.4]
  wire  _T_386; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221306.4]
  wire [26:0] _T_387; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221307.4]
  wire  _T_389; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221309.4]
  wire  sector_hits_0; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221310.4]
  wire  _T_390; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221311.4]
  wire  _T_391; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221312.4]
  wire  _T_392; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221313.4]
  wire [26:0] _T_393; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221314.4]
  wire  _T_395; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221316.4]
  wire  sector_hits_1; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221317.4]
  wire  _T_396; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221318.4]
  wire  _T_397; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221319.4]
  wire  _T_398; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221320.4]
  wire [26:0] _T_399; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221321.4]
  wire  _T_401; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221323.4]
  wire  sector_hits_2; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221324.4]
  wire  _T_402; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221325.4]
  wire  _T_403; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221326.4]
  wire  _T_404; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221327.4]
  wire [26:0] _T_405; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221328.4]
  wire  _T_407; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221330.4]
  wire  sector_hits_3; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221331.4]
  wire  _T_408; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221332.4]
  wire  _T_409; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221333.4]
  wire  _T_410; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221334.4]
  wire [26:0] _T_411; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221335.4]
  wire  _T_413; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221337.4]
  wire  sector_hits_4; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221338.4]
  wire  _T_414; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221339.4]
  wire  _T_415; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221340.4]
  wire  _T_416; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221341.4]
  wire [26:0] _T_417; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221342.4]
  wire  _T_419; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221344.4]
  wire  sector_hits_5; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221345.4]
  wire  _T_420; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221346.4]
  wire  _T_421; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221347.4]
  wire  _T_422; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221348.4]
  wire [26:0] _T_423; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221349.4]
  wire  _T_425; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221351.4]
  wire  sector_hits_6; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221352.4]
  wire  _T_426; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221353.4]
  wire  _T_427; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221354.4]
  wire  _T_428; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221355.4]
  wire [26:0] _T_429; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221356.4]
  wire  _T_431; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221358.4]
  wire  sector_hits_7; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221359.4]
  wire  _T_436; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221364.4]
  wire  _T_438; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221366.4]
  wire  _T_439; // @[TLB.scala 93:28:chipyard.TestHarness.RocketConfig.fir@221367.4]
  wire  _T_443; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221371.4]
  wire  _T_444; // @[TLB.scala 94:40:chipyard.TestHarness.RocketConfig.fir@221372.4]
  wire  superpage_hits_0; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221373.4]
  wire  _T_456; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221385.4]
  wire  _T_458; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221387.4]
  wire  _T_459; // @[TLB.scala 93:28:chipyard.TestHarness.RocketConfig.fir@221388.4]
  wire  _T_463; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221392.4]
  wire  _T_464; // @[TLB.scala 94:40:chipyard.TestHarness.RocketConfig.fir@221393.4]
  wire  superpage_hits_1; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221394.4]
  wire  _T_476; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221406.4]
  wire  _T_478; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221408.4]
  wire  _T_479; // @[TLB.scala 93:28:chipyard.TestHarness.RocketConfig.fir@221409.4]
  wire  _T_483; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221413.4]
  wire  _T_484; // @[TLB.scala 94:40:chipyard.TestHarness.RocketConfig.fir@221414.4]
  wire  superpage_hits_2; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221415.4]
  wire  _T_496; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221427.4]
  wire  _T_498; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221429.4]
  wire  _T_499; // @[TLB.scala 93:28:chipyard.TestHarness.RocketConfig.fir@221430.4]
  wire  _T_503; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221434.4]
  wire  _T_504; // @[TLB.scala 94:40:chipyard.TestHarness.RocketConfig.fir@221435.4]
  wire  superpage_hits_3; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221436.4]
  wire  _GEN_1; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221448.4]
  wire  _GEN_2; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221448.4]
  wire  _GEN_3; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221448.4]
  wire  _T_516; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221448.4]
  wire  hitsVec_0; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221449.4]
  wire  _GEN_5; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221454.4]
  wire  _GEN_6; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221454.4]
  wire  _GEN_7; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221454.4]
  wire  _T_521; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221454.4]
  wire  hitsVec_1; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221455.4]
  wire  _GEN_9; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221460.4]
  wire  _GEN_10; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221460.4]
  wire  _GEN_11; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221460.4]
  wire  _T_526; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221460.4]
  wire  hitsVec_2; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221461.4]
  wire  _GEN_13; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221466.4]
  wire  _GEN_14; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221466.4]
  wire  _GEN_15; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221466.4]
  wire  _T_531; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221466.4]
  wire  hitsVec_3; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221467.4]
  wire  _GEN_17; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221472.4]
  wire  _GEN_18; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221472.4]
  wire  _GEN_19; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221472.4]
  wire  _T_536; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221472.4]
  wire  hitsVec_4; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221473.4]
  wire  _GEN_21; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221478.4]
  wire  _GEN_22; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221478.4]
  wire  _GEN_23; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221478.4]
  wire  _T_541; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221478.4]
  wire  hitsVec_5; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221479.4]
  wire  _GEN_25; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221484.4]
  wire  _GEN_26; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221484.4]
  wire  _GEN_27; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221484.4]
  wire  _T_546; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221484.4]
  wire  hitsVec_6; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221485.4]
  wire  _GEN_29; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221490.4]
  wire  _GEN_30; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221490.4]
  wire  _GEN_31; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221490.4]
  wire  _T_551; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221490.4]
  wire  hitsVec_7; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221491.4]
  wire  hitsVec_8; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221513.4]
  wire  hitsVec_9; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221535.4]
  wire  hitsVec_10; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221557.4]
  wire  hitsVec_11; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221579.4]
  wire  _T_640; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221584.4]
  wire  _T_642; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221586.4]
  wire  _T_647; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221591.4]
  wire  _T_648; // @[TLB.scala 94:40:chipyard.TestHarness.RocketConfig.fir@221592.4]
  wire  _T_649; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221593.4]
  wire  _T_654; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221598.4]
  wire  _T_655; // @[TLB.scala 94:40:chipyard.TestHarness.RocketConfig.fir@221599.4]
  wire  _T_656; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221600.4]
  wire  hitsVec_12; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221601.4]
  wire [5:0] _T_661; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@221606.4]
  wire [12:0] real_hits; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@221613.4]
  wire  _T_668; // @[TLB.scala 211:18:chipyard.TestHarness.RocketConfig.fir@221614.4]
  wire [13:0] hits; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@221615.4]
  wire [33:0] _GEN_33; // @[:chipyard.TestHarness.RocketConfig.fir@221622.4]
  wire [33:0] _GEN_34; // @[:chipyard.TestHarness.RocketConfig.fir@221622.4]
  wire [33:0] _GEN_35; // @[:chipyard.TestHarness.RocketConfig.fir@221622.4]
  wire [33:0] _GEN_37; // @[:chipyard.TestHarness.RocketConfig.fir@221663.4]
  wire [33:0] _GEN_38; // @[:chipyard.TestHarness.RocketConfig.fir@221663.4]
  wire [33:0] _GEN_39; // @[:chipyard.TestHarness.RocketConfig.fir@221663.4]
  wire [33:0] _GEN_41; // @[:chipyard.TestHarness.RocketConfig.fir@221704.4]
  wire [33:0] _GEN_42; // @[:chipyard.TestHarness.RocketConfig.fir@221704.4]
  wire [33:0] _GEN_43; // @[:chipyard.TestHarness.RocketConfig.fir@221704.4]
  wire [33:0] _GEN_45; // @[:chipyard.TestHarness.RocketConfig.fir@221745.4]
  wire [33:0] _GEN_46; // @[:chipyard.TestHarness.RocketConfig.fir@221745.4]
  wire [33:0] _GEN_47; // @[:chipyard.TestHarness.RocketConfig.fir@221745.4]
  wire [33:0] _GEN_49; // @[:chipyard.TestHarness.RocketConfig.fir@221786.4]
  wire [33:0] _GEN_50; // @[:chipyard.TestHarness.RocketConfig.fir@221786.4]
  wire [33:0] _GEN_51; // @[:chipyard.TestHarness.RocketConfig.fir@221786.4]
  wire [33:0] _GEN_53; // @[:chipyard.TestHarness.RocketConfig.fir@221827.4]
  wire [33:0] _GEN_54; // @[:chipyard.TestHarness.RocketConfig.fir@221827.4]
  wire [33:0] _GEN_55; // @[:chipyard.TestHarness.RocketConfig.fir@221827.4]
  wire [33:0] _GEN_57; // @[:chipyard.TestHarness.RocketConfig.fir@221868.4]
  wire [33:0] _GEN_58; // @[:chipyard.TestHarness.RocketConfig.fir@221868.4]
  wire [33:0] _GEN_59; // @[:chipyard.TestHarness.RocketConfig.fir@221868.4]
  wire [33:0] _GEN_61; // @[:chipyard.TestHarness.RocketConfig.fir@221909.4]
  wire [33:0] _GEN_62; // @[:chipyard.TestHarness.RocketConfig.fir@221909.4]
  wire [33:0] _GEN_63; // @[:chipyard.TestHarness.RocketConfig.fir@221909.4]
  wire [26:0] _T_834; // @[TLB.scala 108:28:chipyard.TestHarness.RocketConfig.fir@221988.4]
  wire [26:0] _GEN_952; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@221989.4]
  wire [26:0] _T_835; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@221989.4]
  wire [26:0] _T_841; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@221995.4]
  wire [19:0] _T_843; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@221997.4]
  wire [26:0] _T_864; // @[TLB.scala 108:28:chipyard.TestHarness.RocketConfig.fir@222041.4]
  wire [26:0] _GEN_954; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222042.4]
  wire [26:0] _T_865; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222042.4]
  wire [26:0] _T_871; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222048.4]
  wire [19:0] _T_873; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@222050.4]
  wire [26:0] _T_894; // @[TLB.scala 108:28:chipyard.TestHarness.RocketConfig.fir@222094.4]
  wire [26:0] _GEN_956; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222095.4]
  wire [26:0] _T_895; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222095.4]
  wire [26:0] _T_901; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222101.4]
  wire [19:0] _T_903; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@222103.4]
  wire [26:0] _T_924; // @[TLB.scala 108:28:chipyard.TestHarness.RocketConfig.fir@222147.4]
  wire [26:0] _GEN_958; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222148.4]
  wire [26:0] _T_925; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222148.4]
  wire [26:0] _T_931; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222154.4]
  wire [19:0] _T_933; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@222156.4]
  wire [26:0] _GEN_960; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222201.4]
  wire [26:0] _T_955; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222201.4]
  wire [26:0] _T_961; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222207.4]
  wire [19:0] _T_963; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@222209.4]
  wire [19:0] _T_965; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222211.4]
  wire [19:0] _T_966; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222212.4]
  wire [19:0] _T_967; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222213.4]
  wire [19:0] _T_968; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222214.4]
  wire [19:0] _T_969; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222215.4]
  wire [19:0] _T_970; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222216.4]
  wire [19:0] _T_971; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222217.4]
  wire [19:0] _T_972; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222218.4]
  wire [19:0] _T_973; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222219.4]
  wire [19:0] _T_974; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222220.4]
  wire [19:0] _T_975; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222221.4]
  wire [19:0] _T_976; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222222.4]
  wire [19:0] _T_977; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222223.4]
  wire [19:0] _T_978; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222224.4]
  wire [19:0] _T_979; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222225.4]
  wire [19:0] _T_980; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222226.4]
  wire [19:0] _T_981; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222227.4]
  wire [19:0] _T_982; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222228.4]
  wire [19:0] _T_983; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222229.4]
  wire [19:0] _T_984; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222230.4]
  wire [19:0] _T_985; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222231.4]
  wire [19:0] _T_986; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222232.4]
  wire [19:0] _T_987; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222233.4]
  wire [19:0] _T_988; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222234.4]
  wire [19:0] _T_989; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222235.4]
  wire [19:0] _T_990; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222236.4]
  wire [19:0] ppn; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222237.4]
  wire  _T_992; // @[TLB.scala 215:22:chipyard.TestHarness.RocketConfig.fir@222240.4]
  wire  _T_993; // @[TLB.scala 215:19:chipyard.TestHarness.RocketConfig.fir@222241.4]
  wire  _T_995; // @[TLB.scala 221:25:chipyard.TestHarness.RocketConfig.fir@222248.6]
  wire  _T_996; // @[PTW.scala 69:47:chipyard.TestHarness.RocketConfig.fir@222251.6]
  wire  _T_997; // @[PTW.scala 69:44:chipyard.TestHarness.RocketConfig.fir@222252.6]
  wire  _T_998; // @[PTW.scala 69:38:chipyard.TestHarness.RocketConfig.fir@222253.6]
  wire  _T_999; // @[PTW.scala 69:32:chipyard.TestHarness.RocketConfig.fir@222254.6]
  wire  _T_1000; // @[PTW.scala 69:52:chipyard.TestHarness.RocketConfig.fir@222255.6]
  wire  _T_1001; // @[PTW.scala 73:35:chipyard.TestHarness.RocketConfig.fir@222256.6]
  wire  _T_1007; // @[PTW.scala 74:35:chipyard.TestHarness.RocketConfig.fir@222263.6]
  wire  _T_1008; // @[PTW.scala 74:40:chipyard.TestHarness.RocketConfig.fir@222264.6]
  wire  _T_1014; // @[PTW.scala 75:35:chipyard.TestHarness.RocketConfig.fir@222271.6]
  wire  _T_1015; // @[TLB.scala 234:37:chipyard.TestHarness.RocketConfig.fir@222280.6]
  wire [6:0] _T_1023; // @[TLB.scala 122:24:chipyard.TestHarness.RocketConfig.fir@222292.8]
  wire [33:0] _T_1031; // @[TLB.scala 122:24:chipyard.TestHarness.RocketConfig.fir@222300.8]
  wire  _T_1032; // @[TLB.scala 236:40:chipyard.TestHarness.RocketConfig.fir@222304.8]
  wire  _T_1033; // @[TLB.scala 237:82:chipyard.TestHarness.RocketConfig.fir@222306.10]
  wire  _GEN_66; // @[TLB.scala 237:89:chipyard.TestHarness.RocketConfig.fir@222307.10]
  wire  _T_1049; // @[TLB.scala 237:82:chipyard.TestHarness.RocketConfig.fir@222328.10]
  wire  _GEN_70; // @[TLB.scala 237:89:chipyard.TestHarness.RocketConfig.fir@222329.10]
  wire  _T_1065; // @[TLB.scala 237:82:chipyard.TestHarness.RocketConfig.fir@222350.10]
  wire  _GEN_74; // @[TLB.scala 237:89:chipyard.TestHarness.RocketConfig.fir@222351.10]
  wire  _T_1081; // @[TLB.scala 237:82:chipyard.TestHarness.RocketConfig.fir@222372.10]
  wire  _GEN_78; // @[TLB.scala 237:89:chipyard.TestHarness.RocketConfig.fir@222373.10]
  wire [2:0] _T_1097; // @[TLB.scala 241:22:chipyard.TestHarness.RocketConfig.fir@222396.10]
  wire  _T_1098; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222397.10]
  wire  _T_1099; // @[TLB.scala 243:15:chipyard.TestHarness.RocketConfig.fir@222399.12]
  wire  _GEN_80; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222400.12]
  wire  _GEN_81; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222400.12]
  wire  _GEN_82; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222400.12]
  wire  _GEN_83; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222400.12]
  wire  _GEN_962; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  wire  _GEN_84; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  wire  _GEN_963; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  wire  _GEN_85; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  wire  _GEN_964; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  wire  _GEN_86; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  wire  _GEN_965; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  wire  _GEN_87; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  wire  _GEN_92; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222398.10]
  wire  _GEN_93; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222398.10]
  wire  _GEN_94; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222398.10]
  wire  _GEN_95; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222398.10]
  wire  _T_1115; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222426.10]
  wire  _GEN_102; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222429.12]
  wire  _GEN_103; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222429.12]
  wire  _GEN_104; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222429.12]
  wire  _GEN_105; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222429.12]
  wire  _GEN_106; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222438.12]
  wire  _GEN_107; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222438.12]
  wire  _GEN_108; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222438.12]
  wire  _GEN_109; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222438.12]
  wire  _GEN_114; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222427.10]
  wire  _GEN_115; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222427.10]
  wire  _GEN_116; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222427.10]
  wire  _GEN_117; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222427.10]
  wire  _T_1132; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222455.10]
  wire  _GEN_124; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222458.12]
  wire  _GEN_125; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222458.12]
  wire  _GEN_126; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222458.12]
  wire  _GEN_127; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222458.12]
  wire  _GEN_128; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222467.12]
  wire  _GEN_129; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222467.12]
  wire  _GEN_130; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222467.12]
  wire  _GEN_131; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222467.12]
  wire  _GEN_136; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222456.10]
  wire  _GEN_137; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222456.10]
  wire  _GEN_138; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222456.10]
  wire  _GEN_139; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222456.10]
  wire  _T_1149; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222484.10]
  wire  _GEN_146; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222487.12]
  wire  _GEN_147; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222487.12]
  wire  _GEN_148; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222487.12]
  wire  _GEN_149; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222487.12]
  wire  _GEN_150; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222496.12]
  wire  _GEN_151; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222496.12]
  wire  _GEN_152; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222496.12]
  wire  _GEN_153; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222496.12]
  wire  _GEN_158; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222485.10]
  wire  _GEN_159; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222485.10]
  wire  _GEN_160; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222485.10]
  wire  _GEN_161; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222485.10]
  wire  _T_1166; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222513.10]
  wire  _GEN_168; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222516.12]
  wire  _GEN_169; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222516.12]
  wire  _GEN_170; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222516.12]
  wire  _GEN_171; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222516.12]
  wire  _GEN_172; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222525.12]
  wire  _GEN_173; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222525.12]
  wire  _GEN_174; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222525.12]
  wire  _GEN_175; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222525.12]
  wire  _GEN_180; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222514.10]
  wire  _GEN_181; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222514.10]
  wire  _GEN_182; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222514.10]
  wire  _GEN_183; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222514.10]
  wire  _T_1183; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222542.10]
  wire  _GEN_190; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222545.12]
  wire  _GEN_191; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222545.12]
  wire  _GEN_192; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222545.12]
  wire  _GEN_193; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222545.12]
  wire  _GEN_194; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222554.12]
  wire  _GEN_195; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222554.12]
  wire  _GEN_196; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222554.12]
  wire  _GEN_197; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222554.12]
  wire  _GEN_202; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222543.10]
  wire  _GEN_203; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222543.10]
  wire  _GEN_204; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222543.10]
  wire  _GEN_205; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222543.10]
  wire  _T_1200; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222571.10]
  wire  _GEN_212; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222574.12]
  wire  _GEN_213; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222574.12]
  wire  _GEN_214; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222574.12]
  wire  _GEN_215; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222574.12]
  wire  _GEN_216; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222583.12]
  wire  _GEN_217; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222583.12]
  wire  _GEN_218; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222583.12]
  wire  _GEN_219; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222583.12]
  wire  _GEN_224; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222572.10]
  wire  _GEN_225; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222572.10]
  wire  _GEN_226; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222572.10]
  wire  _GEN_227; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222572.10]
  wire  _T_1217; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222600.10]
  wire  _GEN_234; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222603.12]
  wire  _GEN_235; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222603.12]
  wire  _GEN_236; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222603.12]
  wire  _GEN_237; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222603.12]
  wire  _GEN_238; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222612.12]
  wire  _GEN_239; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222612.12]
  wire  _GEN_240; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222612.12]
  wire  _GEN_241; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222612.12]
  wire  _GEN_246; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222601.10]
  wire  _GEN_247; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222601.10]
  wire  _GEN_248; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222601.10]
  wire  _GEN_249; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222601.10]
  wire  _GEN_258; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_262; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_266; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_270; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_272; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_273; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_274; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_275; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_282; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_283; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_284; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_285; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_292; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_293; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_294; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_295; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_302; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_303; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_304; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_305; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_312; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_313; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_314; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_315; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_322; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_323; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_324; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_325; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_332; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_333; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_334; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_335; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_342; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_343; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_344; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_345; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  wire  _GEN_354; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_358; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_362; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_366; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_370; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_372; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_373; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_374; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_375; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_382; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_383; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_384; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_385; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_392; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_393; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_394; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_395; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_402; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_403; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_404; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_405; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_412; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_413; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_414; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_415; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_422; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_423; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_424; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_425; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_432; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_433; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_434; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_435; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_442; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_443; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_444; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_445; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  wire  _GEN_454; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_458; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_462; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_466; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_470; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_472; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_473; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_474; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_475; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_482; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_483; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_484; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_485; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_492; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_493; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_494; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_495; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_502; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_503; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_504; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_505; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_512; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_513; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_514; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_515; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_522; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_523; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_524; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_525; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_532; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_533; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_534; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_535; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_542; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_543; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_544; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire  _GEN_545; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  wire [5:0] _T_1679; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223651.4]
  wire [13:0] ptw_ae_array; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223659.4]
  wire [5:0] _T_1693; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223666.4]
  wire [12:0] _T_1700; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223673.4]
  wire [12:0] _T_1714; // @[TLB.scala 253:98:chipyard.TestHarness.RocketConfig.fir@223687.4]
  wire [12:0] priv_x_ok; // @[TLB.scala 254:22:chipyard.TestHarness.RocketConfig.fir@223715.4]
  wire [5:0] _T_1757; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223732.4]
  wire [12:0] _T_1764; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223739.4]
  wire [12:0] _T_1793; // @[TLB.scala 257:39:chipyard.TestHarness.RocketConfig.fir@223770.4]
  wire [13:0] x_array; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223771.4]
  wire [13:0] _T_1808; // @[TLB.scala 258:89:chipyard.TestHarness.RocketConfig.fir@223786.4]
  wire [1:0] _T_1825; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@223805.4]
  wire [5:0] _T_1830; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223810.4]
  wire [13:0] _T_1837; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223817.4]
  wire [13:0] px_array; // @[TLB.scala 260:87:chipyard.TestHarness.RocketConfig.fir@223819.4]
  wire [1:0] _T_1853; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@223835.4]
  wire [5:0] _T_1858; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223840.4]
  wire [13:0] c_array; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223847.4]
  wire [39:0] _T_1910; // @[TLB.scala 275:43:chipyard.TestHarness.RocketConfig.fir@223899.4]
  wire  _T_1912; // @[TLB.scala 276:61:chipyard.TestHarness.RocketConfig.fir@223901.4]
  wire  _T_1913; // @[TLB.scala 276:82:chipyard.TestHarness.RocketConfig.fir@223902.4]
  wire  _T_1914; // @[TLB.scala 276:67:chipyard.TestHarness.RocketConfig.fir@223903.4]
  wire  _T_1915; // @[TLB.scala 276:47:chipyard.TestHarness.RocketConfig.fir@223904.4]
  wire  bad_va; // @[TLB.scala 270:117:chipyard.TestHarness.RocketConfig.fir@223906.4]
  wire [13:0] _T_2011; // @[TLB.scala 305:33:chipyard.TestHarness.RocketConfig.fir@224016.4]
  wire [13:0] pf_inst_array; // @[TLB.scala 305:23:chipyard.TestHarness.RocketConfig.fir@224017.4]
  wire  tlb_hit; // @[TLB.scala 307:27:chipyard.TestHarness.RocketConfig.fir@224018.4]
  wire  _T_2012; // @[TLB.scala 308:32:chipyard.TestHarness.RocketConfig.fir@224019.4]
  wire  _T_2013; // @[TLB.scala 308:29:chipyard.TestHarness.RocketConfig.fir@224020.4]
  wire  _T_2014; // @[TLB.scala 308:43:chipyard.TestHarness.RocketConfig.fir@224021.4]
  wire  tlb_miss; // @[TLB.scala 308:40:chipyard.TestHarness.RocketConfig.fir@224022.4]
  reg [6:0] _T_2015; // @[Replacement.scala 42:30:chipyard.TestHarness.RocketConfig.fir@224023.4]
  reg [31:0] _RAND_98;
  reg [2:0] _T_2016; // @[Replacement.scala 42:30:chipyard.TestHarness.RocketConfig.fir@224024.4]
  reg [31:0] _RAND_99;
  wire  _T_2017; // @[TLB.scala 312:22:chipyard.TestHarness.RocketConfig.fir@224025.4]
  wire  _T_2018; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224027.6]
  wire  _T_2019; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224028.6]
  wire  _T_2020; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224029.6]
  wire  _T_2021; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224030.6]
  wire  _T_2022; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224031.6]
  wire  _T_2023; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224032.6]
  wire  _T_2024; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224033.6]
  wire [7:0] _T_2031; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224041.8]
  wire  _T_2034; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@224044.8]
  wire [3:0] _T_2035; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@224045.8]
  wire  _T_2038; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@224048.8]
  wire [1:0] _T_2039; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@224049.8]
  wire [2:0] _T_2042; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224052.8]
  wire [7:0] _T_2043; // @[Replacement.scala 50:28:chipyard.TestHarness.RocketConfig.fir@224053.8]
  wire  _T_2045; // @[Replacement.scala 54:43:chipyard.TestHarness.RocketConfig.fir@224055.8]
  wire [7:0] _T_2047; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224057.8]
  wire [7:0] _T_2048; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224058.8]
  wire [7:0] _T_2049; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224059.8]
  wire [7:0] _T_2050; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224060.8]
  wire [7:0] _T_2051; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224061.8]
  wire [1:0] _T_2052; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224062.8]
  wire  _T_2054; // @[Replacement.scala 54:43:chipyard.TestHarness.RocketConfig.fir@224064.8]
  wire [3:0] _T_2055; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224065.8]
  wire [7:0] _GEN_995; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224066.8]
  wire [7:0] _T_2056; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224066.8]
  wire [7:0] _T_2057; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224067.8]
  wire [7:0] _T_2058; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224068.8]
  wire [7:0] _T_2059; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224069.8]
  wire [7:0] _T_2060; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224070.8]
  wire [2:0] _T_2061; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224071.8]
  wire  _T_2063; // @[Replacement.scala 54:43:chipyard.TestHarness.RocketConfig.fir@224073.8]
  wire [7:0] _T_2064; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224074.8]
  wire [7:0] _T_2065; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224075.8]
  wire [7:0] _T_2066; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224076.8]
  wire [7:0] _T_2067; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224077.8]
  wire [7:0] _T_2068; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224078.8]
  wire [7:0] _T_2069; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224079.8]
  wire  _T_2072; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224084.6]
  wire  _T_2073; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224085.6]
  wire  _T_2074; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224086.6]
  wire [3:0] _T_2077; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224090.8]
  wire  _T_2080; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@224093.8]
  wire [1:0] _T_2081; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@224094.8]
  wire [1:0] _T_2083; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224096.8]
  wire [3:0] _T_2084; // @[Replacement.scala 50:28:chipyard.TestHarness.RocketConfig.fir@224097.8]
  wire  _T_2086; // @[Replacement.scala 54:43:chipyard.TestHarness.RocketConfig.fir@224099.8]
  wire [3:0] _T_2088; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224101.8]
  wire [3:0] _T_2089; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224102.8]
  wire [3:0] _T_2090; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224103.8]
  wire [3:0] _T_2091; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224104.8]
  wire [3:0] _T_2092; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224105.8]
  wire [1:0] _T_2093; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224106.8]
  wire  _T_2095; // @[Replacement.scala 54:43:chipyard.TestHarness.RocketConfig.fir@224108.8]
  wire [3:0] _T_2096; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224109.8]
  wire [3:0] _T_2097; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224110.8]
  wire [3:0] _T_2098; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224111.8]
  wire [3:0] _T_2099; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224112.8]
  wire [3:0] _T_2100; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224113.8]
  wire [3:0] _T_2101; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224114.8]
  wire  _T_2113; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224129.4]
  wire  _T_2115; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224131.4]
  wire  _T_2117; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224133.4]
  wire  _T_2119; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224135.4]
  wire  _T_2120; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224136.4]
  wire  _T_2129; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224145.4]
  wire  _T_2131; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224147.4]
  wire  _T_2133; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224149.4]
  wire  _T_2135; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224151.4]
  wire  _T_2136; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224152.4]
  wire  _T_2137; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224153.4]
  wire  _T_2138; // @[Misc.scala 182:37:chipyard.TestHarness.RocketConfig.fir@224154.4]
  wire  _T_2139; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224155.4]
  wire  _T_2140; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224156.4]
  wire  _T_2150; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224166.4]
  wire  _T_2152; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224168.4]
  wire  _T_2154; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224170.4]
  wire  _T_2156; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224172.4]
  wire  _T_2157; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224173.4]
  wire  _T_2164; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224180.4]
  wire  _T_2166; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224182.4]
  wire  _T_2173; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224189.4]
  wire  _T_2175; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224191.4]
  wire  _T_2177; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224193.4]
  wire  _T_2178; // @[Misc.scala 182:37:chipyard.TestHarness.RocketConfig.fir@224194.4]
  wire  _T_2179; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224195.4]
  wire  _T_2180; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224196.4]
  wire  _T_2181; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224197.4]
  wire  _T_2182; // @[Misc.scala 182:37:chipyard.TestHarness.RocketConfig.fir@224198.4]
  wire  _T_2183; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224199.4]
  wire  _T_2184; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224200.4]
  wire  _T_2186; // @[Misc.scala 182:37:chipyard.TestHarness.RocketConfig.fir@224202.4]
  wire  _T_2187; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224203.4]
  wire  multipleHits; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224204.4]
  wire [13:0] _T_2197; // @[TLB.scala 327:47:chipyard.TestHarness.RocketConfig.fir@224217.4]
  wire  _T_2198; // @[TLB.scala 327:55:chipyard.TestHarness.RocketConfig.fir@224218.4]
  wire [13:0] _T_2204; // @[TLB.scala 330:23:chipyard.TestHarness.RocketConfig.fir@224227.4]
  wire [13:0] _T_2205; // @[TLB.scala 330:33:chipyard.TestHarness.RocketConfig.fir@224228.4]
  wire [13:0] _T_2211; // @[TLB.scala 334:33:chipyard.TestHarness.RocketConfig.fir@224238.4]
  wire  _T_2218; // @[TLB.scala 337:29:chipyard.TestHarness.RocketConfig.fir@224248.4]
  wire  _T_2224; // @[Decoupled.scala 40:37:chipyard.TestHarness.RocketConfig.fir@224259.4]
  wire  _T_2225; // @[TLB.scala 346:25:chipyard.TestHarness.RocketConfig.fir@224260.4]
  wire [3:0] _T_2230; // @[Replacement.scala 65:48:chipyard.TestHarness.RocketConfig.fir@224268.6]
  wire [1:0] _T_2233; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224271.6]
  wire [3:0] _T_2237; // @[Replacement.scala 65:48:chipyard.TestHarness.RocketConfig.fir@224275.6]
  wire [2:0] _T_2240; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224278.6]
  wire [3:0] _T_2244; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224282.6]
  wire  _T_2245; // @[TLB.scala 394:16:chipyard.TestHarness.RocketConfig.fir@224283.6]
  wire [3:0] _T_2246; // @[TLB.scala 394:43:chipyard.TestHarness.RocketConfig.fir@224284.6]
  wire [7:0] _T_2259; // @[Replacement.scala 65:48:chipyard.TestHarness.RocketConfig.fir@224298.6]
  wire [1:0] _T_2262; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224301.6]
  wire [7:0] _T_2266; // @[Replacement.scala 65:48:chipyard.TestHarness.RocketConfig.fir@224305.6]
  wire [2:0] _T_2269; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224308.6]
  wire [7:0] _T_2273; // @[Replacement.scala 65:48:chipyard.TestHarness.RocketConfig.fir@224312.6]
  wire [3:0] _T_2276; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224315.6]
  wire [7:0] _T_2308; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224347.6]
  wire  _T_2309; // @[TLB.scala 394:16:chipyard.TestHarness.RocketConfig.fir@224348.6]
  wire [7:0] _T_2310; // @[TLB.scala 394:43:chipyard.TestHarness.RocketConfig.fir@224349.6]
  wire  _T_2354; // @[TLB.scala 360:17:chipyard.TestHarness.RocketConfig.fir@224408.4]
  wire  _T_2355; // @[TLB.scala 360:28:chipyard.TestHarness.RocketConfig.fir@224409.4]
  wire  _T_2356; // @[TLB.scala 368:14:chipyard.TestHarness.RocketConfig.fir@224417.6]
  wire  _T_2358; // @[TLB.scala 368:72:chipyard.TestHarness.RocketConfig.fir@224419.6]
  wire  _T_2359; // @[TLB.scala 368:34:chipyard.TestHarness.RocketConfig.fir@224420.6]
  wire  _T_2361; // @[TLB.scala 368:13:chipyard.TestHarness.RocketConfig.fir@224422.6]
  wire  _T_2362; // @[TLB.scala 368:13:chipyard.TestHarness.RocketConfig.fir@224423.6]
  wire  _T_2369; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@224438.8]
  wire  _T_2506; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@224736.10]
  wire  _GEN_648; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@224737.10]
  wire  _T_2507; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@224740.10]
  wire  _GEN_649; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@224741.10]
  wire  _T_2508; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@224744.10]
  wire  _GEN_650; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@224745.10]
  wire  _T_2509; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@224748.10]
  wire  _GEN_651; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@224749.10]
  wire  _GEN_652; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224595.8]
  wire  _GEN_653; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224595.8]
  wire  _GEN_654; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224595.8]
  wire  _GEN_655; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224595.8]
  wire  _T_2516; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@224769.8]
  wire  _T_2653; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225067.10]
  wire  _GEN_676; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225068.10]
  wire  _T_2654; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225071.10]
  wire  _GEN_677; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225072.10]
  wire  _T_2655; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225075.10]
  wire  _GEN_678; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225076.10]
  wire  _T_2656; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225079.10]
  wire  _GEN_679; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225080.10]
  wire  _GEN_680; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224926.8]
  wire  _GEN_681; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224926.8]
  wire  _GEN_682; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224926.8]
  wire  _GEN_683; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224926.8]
  wire  _T_2663; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@225100.8]
  wire  _T_2800; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225398.10]
  wire  _GEN_704; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225399.10]
  wire  _T_2801; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225402.10]
  wire  _GEN_705; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225403.10]
  wire  _T_2802; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225406.10]
  wire  _GEN_706; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225407.10]
  wire  _T_2803; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225410.10]
  wire  _GEN_707; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225411.10]
  wire  _GEN_708; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225257.8]
  wire  _GEN_709; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225257.8]
  wire  _GEN_710; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225257.8]
  wire  _GEN_711; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225257.8]
  wire  _T_2810; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@225431.8]
  wire  _T_2947; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225729.10]
  wire  _GEN_732; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225730.10]
  wire  _T_2948; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225733.10]
  wire  _GEN_733; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225734.10]
  wire  _T_2949; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225737.10]
  wire  _GEN_734; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225738.10]
  wire  _T_2950; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225741.10]
  wire  _GEN_735; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225742.10]
  wire  _GEN_736; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225588.8]
  wire  _GEN_737; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225588.8]
  wire  _GEN_738; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225588.8]
  wire  _GEN_739; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225588.8]
  wire  _T_2957; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@225762.8]
  wire  _T_3094; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226060.10]
  wire  _GEN_760; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226061.10]
  wire  _T_3095; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226064.10]
  wire  _GEN_761; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226065.10]
  wire  _T_3096; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226068.10]
  wire  _GEN_762; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226069.10]
  wire  _T_3097; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226072.10]
  wire  _GEN_763; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226073.10]
  wire  _GEN_764; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225919.8]
  wire  _GEN_765; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225919.8]
  wire  _GEN_766; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225919.8]
  wire  _GEN_767; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225919.8]
  wire  _T_3104; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@226093.8]
  wire  _T_3241; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226391.10]
  wire  _GEN_788; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226392.10]
  wire  _T_3242; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226395.10]
  wire  _GEN_789; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226396.10]
  wire  _T_3243; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226399.10]
  wire  _GEN_790; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226400.10]
  wire  _T_3244; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226403.10]
  wire  _GEN_791; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226404.10]
  wire  _GEN_792; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226250.8]
  wire  _GEN_793; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226250.8]
  wire  _GEN_794; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226250.8]
  wire  _GEN_795; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226250.8]
  wire  _T_3251; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@226424.8]
  wire  _T_3388; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226722.10]
  wire  _GEN_816; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226723.10]
  wire  _T_3389; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226726.10]
  wire  _GEN_817; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226727.10]
  wire  _T_3390; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226730.10]
  wire  _GEN_818; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226731.10]
  wire  _T_3391; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226734.10]
  wire  _GEN_819; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226735.10]
  wire  _GEN_820; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226581.8]
  wire  _GEN_821; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226581.8]
  wire  _GEN_822; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226581.8]
  wire  _GEN_823; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226581.8]
  wire  _T_3398; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@226755.8]
  wire  _T_3535; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227053.10]
  wire  _GEN_844; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227054.10]
  wire  _T_3536; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227057.10]
  wire  _GEN_845; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227058.10]
  wire  _T_3537; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227061.10]
  wire  _GEN_846; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227062.10]
  wire  _T_3538; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227065.10]
  wire  _GEN_847; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227066.10]
  wire  _GEN_848; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226912.8]
  wire  _GEN_849; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226912.8]
  wire  _GEN_850; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226912.8]
  wire  _GEN_851; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226912.8]
  wire  _T_3577; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227139.10]
  wire  _GEN_857; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227140.10]
  wire  _GEN_858; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@227103.8]
  wire  _T_3616; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227210.10]
  wire  _GEN_861; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227211.10]
  wire  _GEN_862; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@227174.8]
  wire  _T_3655; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227281.10]
  wire  _GEN_865; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227282.10]
  wire  _GEN_866; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@227245.8]
  wire  _T_3694; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227352.10]
  wire  _GEN_869; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227353.10]
  wire  _GEN_870; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@227316.8]
  wire  _T_3733; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227423.10]
  wire  _GEN_873; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227424.10]
  wire  _GEN_874; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@227387.8]
  wire  _T_3735; // @[TLB.scala 375:24:chipyard.TestHarness.RocketConfig.fir@227433.4]
  package_Anon package_Anon ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@220896.4]
    .io_x_ppn(package_Anon_io_x_ppn),
    .io_x_u(package_Anon_io_x_u),
    .io_x_ae(package_Anon_io_x_ae),
    .io_x_sw(package_Anon_io_x_sw),
    .io_x_sx(package_Anon_io_x_sx),
    .io_x_sr(package_Anon_io_x_sr),
    .io_x_pw(package_Anon_io_x_pw),
    .io_x_px(package_Anon_io_x_px),
    .io_x_pr(package_Anon_io_x_pr),
    .io_x_pal(package_Anon_io_x_pal),
    .io_x_paa(package_Anon_io_x_paa),
    .io_x_eff(package_Anon_io_x_eff),
    .io_x_c(package_Anon_io_x_c),
    .io_y_ppn(package_Anon_io_y_ppn),
    .io_y_u(package_Anon_io_y_u),
    .io_y_ae(package_Anon_io_y_ae),
    .io_y_sw(package_Anon_io_y_sw),
    .io_y_sx(package_Anon_io_y_sx),
    .io_y_sr(package_Anon_io_y_sr),
    .io_y_pw(package_Anon_io_y_pw),
    .io_y_px(package_Anon_io_y_px),
    .io_y_pr(package_Anon_io_y_pr),
    .io_y_pal(package_Anon_io_y_pal),
    .io_y_paa(package_Anon_io_y_paa),
    .io_y_eff(package_Anon_io_y_eff),
    .io_y_c(package_Anon_io_y_c)
  );
  PMPChecker_2 pmp ( // @[TLB.scala 189:19:chipyard.TestHarness.RocketConfig.fir@220923.4]
    .io_prv(pmp_io_prv),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_addr(pmp_io_addr),
    .io_r(pmp_io_r),
    .io_w(pmp_io_w),
    .io_x(pmp_io_x)
  );
  package_Anon package_Anon_1 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221653.4]
    .io_x_ppn(package_Anon_1_io_x_ppn),
    .io_x_u(package_Anon_1_io_x_u),
    .io_x_ae(package_Anon_1_io_x_ae),
    .io_x_sw(package_Anon_1_io_x_sw),
    .io_x_sx(package_Anon_1_io_x_sx),
    .io_x_sr(package_Anon_1_io_x_sr),
    .io_x_pw(package_Anon_1_io_x_pw),
    .io_x_px(package_Anon_1_io_x_px),
    .io_x_pr(package_Anon_1_io_x_pr),
    .io_x_pal(package_Anon_1_io_x_pal),
    .io_x_paa(package_Anon_1_io_x_paa),
    .io_x_eff(package_Anon_1_io_x_eff),
    .io_x_c(package_Anon_1_io_x_c),
    .io_y_ppn(package_Anon_1_io_y_ppn),
    .io_y_u(package_Anon_1_io_y_u),
    .io_y_ae(package_Anon_1_io_y_ae),
    .io_y_sw(package_Anon_1_io_y_sw),
    .io_y_sx(package_Anon_1_io_y_sx),
    .io_y_sr(package_Anon_1_io_y_sr),
    .io_y_pw(package_Anon_1_io_y_pw),
    .io_y_px(package_Anon_1_io_y_px),
    .io_y_pr(package_Anon_1_io_y_pr),
    .io_y_pal(package_Anon_1_io_y_pal),
    .io_y_paa(package_Anon_1_io_y_paa),
    .io_y_eff(package_Anon_1_io_y_eff),
    .io_y_c(package_Anon_1_io_y_c)
  );
  package_Anon package_Anon_2 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221694.4]
    .io_x_ppn(package_Anon_2_io_x_ppn),
    .io_x_u(package_Anon_2_io_x_u),
    .io_x_ae(package_Anon_2_io_x_ae),
    .io_x_sw(package_Anon_2_io_x_sw),
    .io_x_sx(package_Anon_2_io_x_sx),
    .io_x_sr(package_Anon_2_io_x_sr),
    .io_x_pw(package_Anon_2_io_x_pw),
    .io_x_px(package_Anon_2_io_x_px),
    .io_x_pr(package_Anon_2_io_x_pr),
    .io_x_pal(package_Anon_2_io_x_pal),
    .io_x_paa(package_Anon_2_io_x_paa),
    .io_x_eff(package_Anon_2_io_x_eff),
    .io_x_c(package_Anon_2_io_x_c),
    .io_y_ppn(package_Anon_2_io_y_ppn),
    .io_y_u(package_Anon_2_io_y_u),
    .io_y_ae(package_Anon_2_io_y_ae),
    .io_y_sw(package_Anon_2_io_y_sw),
    .io_y_sx(package_Anon_2_io_y_sx),
    .io_y_sr(package_Anon_2_io_y_sr),
    .io_y_pw(package_Anon_2_io_y_pw),
    .io_y_px(package_Anon_2_io_y_px),
    .io_y_pr(package_Anon_2_io_y_pr),
    .io_y_pal(package_Anon_2_io_y_pal),
    .io_y_paa(package_Anon_2_io_y_paa),
    .io_y_eff(package_Anon_2_io_y_eff),
    .io_y_c(package_Anon_2_io_y_c)
  );
  package_Anon package_Anon_3 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221735.4]
    .io_x_ppn(package_Anon_3_io_x_ppn),
    .io_x_u(package_Anon_3_io_x_u),
    .io_x_ae(package_Anon_3_io_x_ae),
    .io_x_sw(package_Anon_3_io_x_sw),
    .io_x_sx(package_Anon_3_io_x_sx),
    .io_x_sr(package_Anon_3_io_x_sr),
    .io_x_pw(package_Anon_3_io_x_pw),
    .io_x_px(package_Anon_3_io_x_px),
    .io_x_pr(package_Anon_3_io_x_pr),
    .io_x_pal(package_Anon_3_io_x_pal),
    .io_x_paa(package_Anon_3_io_x_paa),
    .io_x_eff(package_Anon_3_io_x_eff),
    .io_x_c(package_Anon_3_io_x_c),
    .io_y_ppn(package_Anon_3_io_y_ppn),
    .io_y_u(package_Anon_3_io_y_u),
    .io_y_ae(package_Anon_3_io_y_ae),
    .io_y_sw(package_Anon_3_io_y_sw),
    .io_y_sx(package_Anon_3_io_y_sx),
    .io_y_sr(package_Anon_3_io_y_sr),
    .io_y_pw(package_Anon_3_io_y_pw),
    .io_y_px(package_Anon_3_io_y_px),
    .io_y_pr(package_Anon_3_io_y_pr),
    .io_y_pal(package_Anon_3_io_y_pal),
    .io_y_paa(package_Anon_3_io_y_paa),
    .io_y_eff(package_Anon_3_io_y_eff),
    .io_y_c(package_Anon_3_io_y_c)
  );
  package_Anon package_Anon_4 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221776.4]
    .io_x_ppn(package_Anon_4_io_x_ppn),
    .io_x_u(package_Anon_4_io_x_u),
    .io_x_ae(package_Anon_4_io_x_ae),
    .io_x_sw(package_Anon_4_io_x_sw),
    .io_x_sx(package_Anon_4_io_x_sx),
    .io_x_sr(package_Anon_4_io_x_sr),
    .io_x_pw(package_Anon_4_io_x_pw),
    .io_x_px(package_Anon_4_io_x_px),
    .io_x_pr(package_Anon_4_io_x_pr),
    .io_x_pal(package_Anon_4_io_x_pal),
    .io_x_paa(package_Anon_4_io_x_paa),
    .io_x_eff(package_Anon_4_io_x_eff),
    .io_x_c(package_Anon_4_io_x_c),
    .io_y_ppn(package_Anon_4_io_y_ppn),
    .io_y_u(package_Anon_4_io_y_u),
    .io_y_ae(package_Anon_4_io_y_ae),
    .io_y_sw(package_Anon_4_io_y_sw),
    .io_y_sx(package_Anon_4_io_y_sx),
    .io_y_sr(package_Anon_4_io_y_sr),
    .io_y_pw(package_Anon_4_io_y_pw),
    .io_y_px(package_Anon_4_io_y_px),
    .io_y_pr(package_Anon_4_io_y_pr),
    .io_y_pal(package_Anon_4_io_y_pal),
    .io_y_paa(package_Anon_4_io_y_paa),
    .io_y_eff(package_Anon_4_io_y_eff),
    .io_y_c(package_Anon_4_io_y_c)
  );
  package_Anon package_Anon_5 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221817.4]
    .io_x_ppn(package_Anon_5_io_x_ppn),
    .io_x_u(package_Anon_5_io_x_u),
    .io_x_ae(package_Anon_5_io_x_ae),
    .io_x_sw(package_Anon_5_io_x_sw),
    .io_x_sx(package_Anon_5_io_x_sx),
    .io_x_sr(package_Anon_5_io_x_sr),
    .io_x_pw(package_Anon_5_io_x_pw),
    .io_x_px(package_Anon_5_io_x_px),
    .io_x_pr(package_Anon_5_io_x_pr),
    .io_x_pal(package_Anon_5_io_x_pal),
    .io_x_paa(package_Anon_5_io_x_paa),
    .io_x_eff(package_Anon_5_io_x_eff),
    .io_x_c(package_Anon_5_io_x_c),
    .io_y_ppn(package_Anon_5_io_y_ppn),
    .io_y_u(package_Anon_5_io_y_u),
    .io_y_ae(package_Anon_5_io_y_ae),
    .io_y_sw(package_Anon_5_io_y_sw),
    .io_y_sx(package_Anon_5_io_y_sx),
    .io_y_sr(package_Anon_5_io_y_sr),
    .io_y_pw(package_Anon_5_io_y_pw),
    .io_y_px(package_Anon_5_io_y_px),
    .io_y_pr(package_Anon_5_io_y_pr),
    .io_y_pal(package_Anon_5_io_y_pal),
    .io_y_paa(package_Anon_5_io_y_paa),
    .io_y_eff(package_Anon_5_io_y_eff),
    .io_y_c(package_Anon_5_io_y_c)
  );
  package_Anon package_Anon_6 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221858.4]
    .io_x_ppn(package_Anon_6_io_x_ppn),
    .io_x_u(package_Anon_6_io_x_u),
    .io_x_ae(package_Anon_6_io_x_ae),
    .io_x_sw(package_Anon_6_io_x_sw),
    .io_x_sx(package_Anon_6_io_x_sx),
    .io_x_sr(package_Anon_6_io_x_sr),
    .io_x_pw(package_Anon_6_io_x_pw),
    .io_x_px(package_Anon_6_io_x_px),
    .io_x_pr(package_Anon_6_io_x_pr),
    .io_x_pal(package_Anon_6_io_x_pal),
    .io_x_paa(package_Anon_6_io_x_paa),
    .io_x_eff(package_Anon_6_io_x_eff),
    .io_x_c(package_Anon_6_io_x_c),
    .io_y_ppn(package_Anon_6_io_y_ppn),
    .io_y_u(package_Anon_6_io_y_u),
    .io_y_ae(package_Anon_6_io_y_ae),
    .io_y_sw(package_Anon_6_io_y_sw),
    .io_y_sx(package_Anon_6_io_y_sx),
    .io_y_sr(package_Anon_6_io_y_sr),
    .io_y_pw(package_Anon_6_io_y_pw),
    .io_y_px(package_Anon_6_io_y_px),
    .io_y_pr(package_Anon_6_io_y_pr),
    .io_y_pal(package_Anon_6_io_y_pal),
    .io_y_paa(package_Anon_6_io_y_paa),
    .io_y_eff(package_Anon_6_io_y_eff),
    .io_y_c(package_Anon_6_io_y_c)
  );
  package_Anon package_Anon_7 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221899.4]
    .io_x_ppn(package_Anon_7_io_x_ppn),
    .io_x_u(package_Anon_7_io_x_u),
    .io_x_ae(package_Anon_7_io_x_ae),
    .io_x_sw(package_Anon_7_io_x_sw),
    .io_x_sx(package_Anon_7_io_x_sx),
    .io_x_sr(package_Anon_7_io_x_sr),
    .io_x_pw(package_Anon_7_io_x_pw),
    .io_x_px(package_Anon_7_io_x_px),
    .io_x_pr(package_Anon_7_io_x_pr),
    .io_x_pal(package_Anon_7_io_x_pal),
    .io_x_paa(package_Anon_7_io_x_paa),
    .io_x_eff(package_Anon_7_io_x_eff),
    .io_x_c(package_Anon_7_io_x_c),
    .io_y_ppn(package_Anon_7_io_y_ppn),
    .io_y_u(package_Anon_7_io_y_u),
    .io_y_ae(package_Anon_7_io_y_ae),
    .io_y_sw(package_Anon_7_io_y_sw),
    .io_y_sx(package_Anon_7_io_y_sx),
    .io_y_sr(package_Anon_7_io_y_sr),
    .io_y_pw(package_Anon_7_io_y_pw),
    .io_y_px(package_Anon_7_io_y_px),
    .io_y_pr(package_Anon_7_io_y_pr),
    .io_y_pal(package_Anon_7_io_y_pal),
    .io_y_paa(package_Anon_7_io_y_paa),
    .io_y_eff(package_Anon_7_io_y_eff),
    .io_y_c(package_Anon_7_io_y_c)
  );
  package_Anon package_Anon_8 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221940.4]
    .io_x_ppn(package_Anon_8_io_x_ppn),
    .io_x_u(package_Anon_8_io_x_u),
    .io_x_ae(package_Anon_8_io_x_ae),
    .io_x_sw(package_Anon_8_io_x_sw),
    .io_x_sx(package_Anon_8_io_x_sx),
    .io_x_sr(package_Anon_8_io_x_sr),
    .io_x_pw(package_Anon_8_io_x_pw),
    .io_x_px(package_Anon_8_io_x_px),
    .io_x_pr(package_Anon_8_io_x_pr),
    .io_x_pal(package_Anon_8_io_x_pal),
    .io_x_paa(package_Anon_8_io_x_paa),
    .io_x_eff(package_Anon_8_io_x_eff),
    .io_x_c(package_Anon_8_io_x_c),
    .io_y_ppn(package_Anon_8_io_y_ppn),
    .io_y_u(package_Anon_8_io_y_u),
    .io_y_ae(package_Anon_8_io_y_ae),
    .io_y_sw(package_Anon_8_io_y_sw),
    .io_y_sx(package_Anon_8_io_y_sx),
    .io_y_sr(package_Anon_8_io_y_sr),
    .io_y_pw(package_Anon_8_io_y_pw),
    .io_y_px(package_Anon_8_io_y_px),
    .io_y_pr(package_Anon_8_io_y_pr),
    .io_y_pal(package_Anon_8_io_y_pal),
    .io_y_paa(package_Anon_8_io_y_paa),
    .io_y_eff(package_Anon_8_io_y_eff),
    .io_y_c(package_Anon_8_io_y_c)
  );
  package_Anon package_Anon_9 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@221980.4]
    .io_x_ppn(package_Anon_9_io_x_ppn),
    .io_x_u(package_Anon_9_io_x_u),
    .io_x_ae(package_Anon_9_io_x_ae),
    .io_x_sw(package_Anon_9_io_x_sw),
    .io_x_sx(package_Anon_9_io_x_sx),
    .io_x_sr(package_Anon_9_io_x_sr),
    .io_x_pw(package_Anon_9_io_x_pw),
    .io_x_px(package_Anon_9_io_x_px),
    .io_x_pr(package_Anon_9_io_x_pr),
    .io_x_pal(package_Anon_9_io_x_pal),
    .io_x_paa(package_Anon_9_io_x_paa),
    .io_x_eff(package_Anon_9_io_x_eff),
    .io_x_c(package_Anon_9_io_x_c),
    .io_y_ppn(package_Anon_9_io_y_ppn),
    .io_y_u(package_Anon_9_io_y_u),
    .io_y_ae(package_Anon_9_io_y_ae),
    .io_y_sw(package_Anon_9_io_y_sw),
    .io_y_sx(package_Anon_9_io_y_sx),
    .io_y_sr(package_Anon_9_io_y_sr),
    .io_y_pw(package_Anon_9_io_y_pw),
    .io_y_px(package_Anon_9_io_y_px),
    .io_y_pr(package_Anon_9_io_y_pr),
    .io_y_pal(package_Anon_9_io_y_pal),
    .io_y_paa(package_Anon_9_io_y_paa),
    .io_y_eff(package_Anon_9_io_y_eff),
    .io_y_c(package_Anon_9_io_y_c)
  );
  package_Anon package_Anon_10 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222033.4]
    .io_x_ppn(package_Anon_10_io_x_ppn),
    .io_x_u(package_Anon_10_io_x_u),
    .io_x_ae(package_Anon_10_io_x_ae),
    .io_x_sw(package_Anon_10_io_x_sw),
    .io_x_sx(package_Anon_10_io_x_sx),
    .io_x_sr(package_Anon_10_io_x_sr),
    .io_x_pw(package_Anon_10_io_x_pw),
    .io_x_px(package_Anon_10_io_x_px),
    .io_x_pr(package_Anon_10_io_x_pr),
    .io_x_pal(package_Anon_10_io_x_pal),
    .io_x_paa(package_Anon_10_io_x_paa),
    .io_x_eff(package_Anon_10_io_x_eff),
    .io_x_c(package_Anon_10_io_x_c),
    .io_y_ppn(package_Anon_10_io_y_ppn),
    .io_y_u(package_Anon_10_io_y_u),
    .io_y_ae(package_Anon_10_io_y_ae),
    .io_y_sw(package_Anon_10_io_y_sw),
    .io_y_sx(package_Anon_10_io_y_sx),
    .io_y_sr(package_Anon_10_io_y_sr),
    .io_y_pw(package_Anon_10_io_y_pw),
    .io_y_px(package_Anon_10_io_y_px),
    .io_y_pr(package_Anon_10_io_y_pr),
    .io_y_pal(package_Anon_10_io_y_pal),
    .io_y_paa(package_Anon_10_io_y_paa),
    .io_y_eff(package_Anon_10_io_y_eff),
    .io_y_c(package_Anon_10_io_y_c)
  );
  package_Anon package_Anon_11 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222086.4]
    .io_x_ppn(package_Anon_11_io_x_ppn),
    .io_x_u(package_Anon_11_io_x_u),
    .io_x_ae(package_Anon_11_io_x_ae),
    .io_x_sw(package_Anon_11_io_x_sw),
    .io_x_sx(package_Anon_11_io_x_sx),
    .io_x_sr(package_Anon_11_io_x_sr),
    .io_x_pw(package_Anon_11_io_x_pw),
    .io_x_px(package_Anon_11_io_x_px),
    .io_x_pr(package_Anon_11_io_x_pr),
    .io_x_pal(package_Anon_11_io_x_pal),
    .io_x_paa(package_Anon_11_io_x_paa),
    .io_x_eff(package_Anon_11_io_x_eff),
    .io_x_c(package_Anon_11_io_x_c),
    .io_y_ppn(package_Anon_11_io_y_ppn),
    .io_y_u(package_Anon_11_io_y_u),
    .io_y_ae(package_Anon_11_io_y_ae),
    .io_y_sw(package_Anon_11_io_y_sw),
    .io_y_sx(package_Anon_11_io_y_sx),
    .io_y_sr(package_Anon_11_io_y_sr),
    .io_y_pw(package_Anon_11_io_y_pw),
    .io_y_px(package_Anon_11_io_y_px),
    .io_y_pr(package_Anon_11_io_y_pr),
    .io_y_pal(package_Anon_11_io_y_pal),
    .io_y_paa(package_Anon_11_io_y_paa),
    .io_y_eff(package_Anon_11_io_y_eff),
    .io_y_c(package_Anon_11_io_y_c)
  );
  package_Anon package_Anon_12 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222139.4]
    .io_x_ppn(package_Anon_12_io_x_ppn),
    .io_x_u(package_Anon_12_io_x_u),
    .io_x_ae(package_Anon_12_io_x_ae),
    .io_x_sw(package_Anon_12_io_x_sw),
    .io_x_sx(package_Anon_12_io_x_sx),
    .io_x_sr(package_Anon_12_io_x_sr),
    .io_x_pw(package_Anon_12_io_x_pw),
    .io_x_px(package_Anon_12_io_x_px),
    .io_x_pr(package_Anon_12_io_x_pr),
    .io_x_pal(package_Anon_12_io_x_pal),
    .io_x_paa(package_Anon_12_io_x_paa),
    .io_x_eff(package_Anon_12_io_x_eff),
    .io_x_c(package_Anon_12_io_x_c),
    .io_y_ppn(package_Anon_12_io_y_ppn),
    .io_y_u(package_Anon_12_io_y_u),
    .io_y_ae(package_Anon_12_io_y_ae),
    .io_y_sw(package_Anon_12_io_y_sw),
    .io_y_sx(package_Anon_12_io_y_sx),
    .io_y_sr(package_Anon_12_io_y_sr),
    .io_y_pw(package_Anon_12_io_y_pw),
    .io_y_px(package_Anon_12_io_y_px),
    .io_y_pr(package_Anon_12_io_y_pr),
    .io_y_pal(package_Anon_12_io_y_pal),
    .io_y_paa(package_Anon_12_io_y_paa),
    .io_y_eff(package_Anon_12_io_y_eff),
    .io_y_c(package_Anon_12_io_y_c)
  );
  package_Anon package_Anon_13 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222192.4]
    .io_x_ppn(package_Anon_13_io_x_ppn),
    .io_x_u(package_Anon_13_io_x_u),
    .io_x_ae(package_Anon_13_io_x_ae),
    .io_x_sw(package_Anon_13_io_x_sw),
    .io_x_sx(package_Anon_13_io_x_sx),
    .io_x_sr(package_Anon_13_io_x_sr),
    .io_x_pw(package_Anon_13_io_x_pw),
    .io_x_px(package_Anon_13_io_x_px),
    .io_x_pr(package_Anon_13_io_x_pr),
    .io_x_pal(package_Anon_13_io_x_pal),
    .io_x_paa(package_Anon_13_io_x_paa),
    .io_x_eff(package_Anon_13_io_x_eff),
    .io_x_c(package_Anon_13_io_x_c),
    .io_y_ppn(package_Anon_13_io_y_ppn),
    .io_y_u(package_Anon_13_io_y_u),
    .io_y_ae(package_Anon_13_io_y_ae),
    .io_y_sw(package_Anon_13_io_y_sw),
    .io_y_sx(package_Anon_13_io_y_sx),
    .io_y_sr(package_Anon_13_io_y_sr),
    .io_y_pw(package_Anon_13_io_y_pw),
    .io_y_px(package_Anon_13_io_y_px),
    .io_y_pr(package_Anon_13_io_y_pr),
    .io_y_pal(package_Anon_13_io_y_pal),
    .io_y_paa(package_Anon_13_io_y_paa),
    .io_y_eff(package_Anon_13_io_y_eff),
    .io_y_c(package_Anon_13_io_y_c)
  );
  package_Anon package_Anon_14 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222667.4]
    .io_x_ppn(package_Anon_14_io_x_ppn),
    .io_x_u(package_Anon_14_io_x_u),
    .io_x_ae(package_Anon_14_io_x_ae),
    .io_x_sw(package_Anon_14_io_x_sw),
    .io_x_sx(package_Anon_14_io_x_sx),
    .io_x_sr(package_Anon_14_io_x_sr),
    .io_x_pw(package_Anon_14_io_x_pw),
    .io_x_px(package_Anon_14_io_x_px),
    .io_x_pr(package_Anon_14_io_x_pr),
    .io_x_pal(package_Anon_14_io_x_pal),
    .io_x_paa(package_Anon_14_io_x_paa),
    .io_x_eff(package_Anon_14_io_x_eff),
    .io_x_c(package_Anon_14_io_x_c),
    .io_y_ppn(package_Anon_14_io_y_ppn),
    .io_y_u(package_Anon_14_io_y_u),
    .io_y_ae(package_Anon_14_io_y_ae),
    .io_y_sw(package_Anon_14_io_y_sw),
    .io_y_sx(package_Anon_14_io_y_sx),
    .io_y_sr(package_Anon_14_io_y_sr),
    .io_y_pw(package_Anon_14_io_y_pw),
    .io_y_px(package_Anon_14_io_y_px),
    .io_y_pr(package_Anon_14_io_y_pr),
    .io_y_pal(package_Anon_14_io_y_pal),
    .io_y_paa(package_Anon_14_io_y_paa),
    .io_y_eff(package_Anon_14_io_y_eff),
    .io_y_c(package_Anon_14_io_y_c)
  );
  package_Anon package_Anon_15 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222708.4]
    .io_x_ppn(package_Anon_15_io_x_ppn),
    .io_x_u(package_Anon_15_io_x_u),
    .io_x_ae(package_Anon_15_io_x_ae),
    .io_x_sw(package_Anon_15_io_x_sw),
    .io_x_sx(package_Anon_15_io_x_sx),
    .io_x_sr(package_Anon_15_io_x_sr),
    .io_x_pw(package_Anon_15_io_x_pw),
    .io_x_px(package_Anon_15_io_x_px),
    .io_x_pr(package_Anon_15_io_x_pr),
    .io_x_pal(package_Anon_15_io_x_pal),
    .io_x_paa(package_Anon_15_io_x_paa),
    .io_x_eff(package_Anon_15_io_x_eff),
    .io_x_c(package_Anon_15_io_x_c),
    .io_y_ppn(package_Anon_15_io_y_ppn),
    .io_y_u(package_Anon_15_io_y_u),
    .io_y_ae(package_Anon_15_io_y_ae),
    .io_y_sw(package_Anon_15_io_y_sw),
    .io_y_sx(package_Anon_15_io_y_sx),
    .io_y_sr(package_Anon_15_io_y_sr),
    .io_y_pw(package_Anon_15_io_y_pw),
    .io_y_px(package_Anon_15_io_y_px),
    .io_y_pr(package_Anon_15_io_y_pr),
    .io_y_pal(package_Anon_15_io_y_pal),
    .io_y_paa(package_Anon_15_io_y_paa),
    .io_y_eff(package_Anon_15_io_y_eff),
    .io_y_c(package_Anon_15_io_y_c)
  );
  package_Anon package_Anon_16 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222749.4]
    .io_x_ppn(package_Anon_16_io_x_ppn),
    .io_x_u(package_Anon_16_io_x_u),
    .io_x_ae(package_Anon_16_io_x_ae),
    .io_x_sw(package_Anon_16_io_x_sw),
    .io_x_sx(package_Anon_16_io_x_sx),
    .io_x_sr(package_Anon_16_io_x_sr),
    .io_x_pw(package_Anon_16_io_x_pw),
    .io_x_px(package_Anon_16_io_x_px),
    .io_x_pr(package_Anon_16_io_x_pr),
    .io_x_pal(package_Anon_16_io_x_pal),
    .io_x_paa(package_Anon_16_io_x_paa),
    .io_x_eff(package_Anon_16_io_x_eff),
    .io_x_c(package_Anon_16_io_x_c),
    .io_y_ppn(package_Anon_16_io_y_ppn),
    .io_y_u(package_Anon_16_io_y_u),
    .io_y_ae(package_Anon_16_io_y_ae),
    .io_y_sw(package_Anon_16_io_y_sw),
    .io_y_sx(package_Anon_16_io_y_sx),
    .io_y_sr(package_Anon_16_io_y_sr),
    .io_y_pw(package_Anon_16_io_y_pw),
    .io_y_px(package_Anon_16_io_y_px),
    .io_y_pr(package_Anon_16_io_y_pr),
    .io_y_pal(package_Anon_16_io_y_pal),
    .io_y_paa(package_Anon_16_io_y_paa),
    .io_y_eff(package_Anon_16_io_y_eff),
    .io_y_c(package_Anon_16_io_y_c)
  );
  package_Anon package_Anon_17 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222790.4]
    .io_x_ppn(package_Anon_17_io_x_ppn),
    .io_x_u(package_Anon_17_io_x_u),
    .io_x_ae(package_Anon_17_io_x_ae),
    .io_x_sw(package_Anon_17_io_x_sw),
    .io_x_sx(package_Anon_17_io_x_sx),
    .io_x_sr(package_Anon_17_io_x_sr),
    .io_x_pw(package_Anon_17_io_x_pw),
    .io_x_px(package_Anon_17_io_x_px),
    .io_x_pr(package_Anon_17_io_x_pr),
    .io_x_pal(package_Anon_17_io_x_pal),
    .io_x_paa(package_Anon_17_io_x_paa),
    .io_x_eff(package_Anon_17_io_x_eff),
    .io_x_c(package_Anon_17_io_x_c),
    .io_y_ppn(package_Anon_17_io_y_ppn),
    .io_y_u(package_Anon_17_io_y_u),
    .io_y_ae(package_Anon_17_io_y_ae),
    .io_y_sw(package_Anon_17_io_y_sw),
    .io_y_sx(package_Anon_17_io_y_sx),
    .io_y_sr(package_Anon_17_io_y_sr),
    .io_y_pw(package_Anon_17_io_y_pw),
    .io_y_px(package_Anon_17_io_y_px),
    .io_y_pr(package_Anon_17_io_y_pr),
    .io_y_pal(package_Anon_17_io_y_pal),
    .io_y_paa(package_Anon_17_io_y_paa),
    .io_y_eff(package_Anon_17_io_y_eff),
    .io_y_c(package_Anon_17_io_y_c)
  );
  package_Anon package_Anon_18 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222831.4]
    .io_x_ppn(package_Anon_18_io_x_ppn),
    .io_x_u(package_Anon_18_io_x_u),
    .io_x_ae(package_Anon_18_io_x_ae),
    .io_x_sw(package_Anon_18_io_x_sw),
    .io_x_sx(package_Anon_18_io_x_sx),
    .io_x_sr(package_Anon_18_io_x_sr),
    .io_x_pw(package_Anon_18_io_x_pw),
    .io_x_px(package_Anon_18_io_x_px),
    .io_x_pr(package_Anon_18_io_x_pr),
    .io_x_pal(package_Anon_18_io_x_pal),
    .io_x_paa(package_Anon_18_io_x_paa),
    .io_x_eff(package_Anon_18_io_x_eff),
    .io_x_c(package_Anon_18_io_x_c),
    .io_y_ppn(package_Anon_18_io_y_ppn),
    .io_y_u(package_Anon_18_io_y_u),
    .io_y_ae(package_Anon_18_io_y_ae),
    .io_y_sw(package_Anon_18_io_y_sw),
    .io_y_sx(package_Anon_18_io_y_sx),
    .io_y_sr(package_Anon_18_io_y_sr),
    .io_y_pw(package_Anon_18_io_y_pw),
    .io_y_px(package_Anon_18_io_y_px),
    .io_y_pr(package_Anon_18_io_y_pr),
    .io_y_pal(package_Anon_18_io_y_pal),
    .io_y_paa(package_Anon_18_io_y_paa),
    .io_y_eff(package_Anon_18_io_y_eff),
    .io_y_c(package_Anon_18_io_y_c)
  );
  package_Anon package_Anon_19 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222872.4]
    .io_x_ppn(package_Anon_19_io_x_ppn),
    .io_x_u(package_Anon_19_io_x_u),
    .io_x_ae(package_Anon_19_io_x_ae),
    .io_x_sw(package_Anon_19_io_x_sw),
    .io_x_sx(package_Anon_19_io_x_sx),
    .io_x_sr(package_Anon_19_io_x_sr),
    .io_x_pw(package_Anon_19_io_x_pw),
    .io_x_px(package_Anon_19_io_x_px),
    .io_x_pr(package_Anon_19_io_x_pr),
    .io_x_pal(package_Anon_19_io_x_pal),
    .io_x_paa(package_Anon_19_io_x_paa),
    .io_x_eff(package_Anon_19_io_x_eff),
    .io_x_c(package_Anon_19_io_x_c),
    .io_y_ppn(package_Anon_19_io_y_ppn),
    .io_y_u(package_Anon_19_io_y_u),
    .io_y_ae(package_Anon_19_io_y_ae),
    .io_y_sw(package_Anon_19_io_y_sw),
    .io_y_sx(package_Anon_19_io_y_sx),
    .io_y_sr(package_Anon_19_io_y_sr),
    .io_y_pw(package_Anon_19_io_y_pw),
    .io_y_px(package_Anon_19_io_y_px),
    .io_y_pr(package_Anon_19_io_y_pr),
    .io_y_pal(package_Anon_19_io_y_pal),
    .io_y_paa(package_Anon_19_io_y_paa),
    .io_y_eff(package_Anon_19_io_y_eff),
    .io_y_c(package_Anon_19_io_y_c)
  );
  package_Anon package_Anon_20 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222913.4]
    .io_x_ppn(package_Anon_20_io_x_ppn),
    .io_x_u(package_Anon_20_io_x_u),
    .io_x_ae(package_Anon_20_io_x_ae),
    .io_x_sw(package_Anon_20_io_x_sw),
    .io_x_sx(package_Anon_20_io_x_sx),
    .io_x_sr(package_Anon_20_io_x_sr),
    .io_x_pw(package_Anon_20_io_x_pw),
    .io_x_px(package_Anon_20_io_x_px),
    .io_x_pr(package_Anon_20_io_x_pr),
    .io_x_pal(package_Anon_20_io_x_pal),
    .io_x_paa(package_Anon_20_io_x_paa),
    .io_x_eff(package_Anon_20_io_x_eff),
    .io_x_c(package_Anon_20_io_x_c),
    .io_y_ppn(package_Anon_20_io_y_ppn),
    .io_y_u(package_Anon_20_io_y_u),
    .io_y_ae(package_Anon_20_io_y_ae),
    .io_y_sw(package_Anon_20_io_y_sw),
    .io_y_sx(package_Anon_20_io_y_sx),
    .io_y_sr(package_Anon_20_io_y_sr),
    .io_y_pw(package_Anon_20_io_y_pw),
    .io_y_px(package_Anon_20_io_y_px),
    .io_y_pr(package_Anon_20_io_y_pr),
    .io_y_pal(package_Anon_20_io_y_pal),
    .io_y_paa(package_Anon_20_io_y_paa),
    .io_y_eff(package_Anon_20_io_y_eff),
    .io_y_c(package_Anon_20_io_y_c)
  );
  package_Anon package_Anon_21 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222954.4]
    .io_x_ppn(package_Anon_21_io_x_ppn),
    .io_x_u(package_Anon_21_io_x_u),
    .io_x_ae(package_Anon_21_io_x_ae),
    .io_x_sw(package_Anon_21_io_x_sw),
    .io_x_sx(package_Anon_21_io_x_sx),
    .io_x_sr(package_Anon_21_io_x_sr),
    .io_x_pw(package_Anon_21_io_x_pw),
    .io_x_px(package_Anon_21_io_x_px),
    .io_x_pr(package_Anon_21_io_x_pr),
    .io_x_pal(package_Anon_21_io_x_pal),
    .io_x_paa(package_Anon_21_io_x_paa),
    .io_x_eff(package_Anon_21_io_x_eff),
    .io_x_c(package_Anon_21_io_x_c),
    .io_y_ppn(package_Anon_21_io_y_ppn),
    .io_y_u(package_Anon_21_io_y_u),
    .io_y_ae(package_Anon_21_io_y_ae),
    .io_y_sw(package_Anon_21_io_y_sw),
    .io_y_sx(package_Anon_21_io_y_sx),
    .io_y_sr(package_Anon_21_io_y_sr),
    .io_y_pw(package_Anon_21_io_y_pw),
    .io_y_px(package_Anon_21_io_y_px),
    .io_y_pr(package_Anon_21_io_y_pr),
    .io_y_pal(package_Anon_21_io_y_pal),
    .io_y_paa(package_Anon_21_io_y_paa),
    .io_y_eff(package_Anon_21_io_y_eff),
    .io_y_c(package_Anon_21_io_y_c)
  );
  package_Anon package_Anon_22 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@222994.4]
    .io_x_ppn(package_Anon_22_io_x_ppn),
    .io_x_u(package_Anon_22_io_x_u),
    .io_x_ae(package_Anon_22_io_x_ae),
    .io_x_sw(package_Anon_22_io_x_sw),
    .io_x_sx(package_Anon_22_io_x_sx),
    .io_x_sr(package_Anon_22_io_x_sr),
    .io_x_pw(package_Anon_22_io_x_pw),
    .io_x_px(package_Anon_22_io_x_px),
    .io_x_pr(package_Anon_22_io_x_pr),
    .io_x_pal(package_Anon_22_io_x_pal),
    .io_x_paa(package_Anon_22_io_x_paa),
    .io_x_eff(package_Anon_22_io_x_eff),
    .io_x_c(package_Anon_22_io_x_c),
    .io_y_ppn(package_Anon_22_io_y_ppn),
    .io_y_u(package_Anon_22_io_y_u),
    .io_y_ae(package_Anon_22_io_y_ae),
    .io_y_sw(package_Anon_22_io_y_sw),
    .io_y_sx(package_Anon_22_io_y_sx),
    .io_y_sr(package_Anon_22_io_y_sr),
    .io_y_pw(package_Anon_22_io_y_pw),
    .io_y_px(package_Anon_22_io_y_px),
    .io_y_pr(package_Anon_22_io_y_pr),
    .io_y_pal(package_Anon_22_io_y_pal),
    .io_y_paa(package_Anon_22_io_y_paa),
    .io_y_eff(package_Anon_22_io_y_eff),
    .io_y_c(package_Anon_22_io_y_c)
  );
  package_Anon package_Anon_23 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223034.4]
    .io_x_ppn(package_Anon_23_io_x_ppn),
    .io_x_u(package_Anon_23_io_x_u),
    .io_x_ae(package_Anon_23_io_x_ae),
    .io_x_sw(package_Anon_23_io_x_sw),
    .io_x_sx(package_Anon_23_io_x_sx),
    .io_x_sr(package_Anon_23_io_x_sr),
    .io_x_pw(package_Anon_23_io_x_pw),
    .io_x_px(package_Anon_23_io_x_px),
    .io_x_pr(package_Anon_23_io_x_pr),
    .io_x_pal(package_Anon_23_io_x_pal),
    .io_x_paa(package_Anon_23_io_x_paa),
    .io_x_eff(package_Anon_23_io_x_eff),
    .io_x_c(package_Anon_23_io_x_c),
    .io_y_ppn(package_Anon_23_io_y_ppn),
    .io_y_u(package_Anon_23_io_y_u),
    .io_y_ae(package_Anon_23_io_y_ae),
    .io_y_sw(package_Anon_23_io_y_sw),
    .io_y_sx(package_Anon_23_io_y_sx),
    .io_y_sr(package_Anon_23_io_y_sr),
    .io_y_pw(package_Anon_23_io_y_pw),
    .io_y_px(package_Anon_23_io_y_px),
    .io_y_pr(package_Anon_23_io_y_pr),
    .io_y_pal(package_Anon_23_io_y_pal),
    .io_y_paa(package_Anon_23_io_y_paa),
    .io_y_eff(package_Anon_23_io_y_eff),
    .io_y_c(package_Anon_23_io_y_c)
  );
  package_Anon package_Anon_24 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223074.4]
    .io_x_ppn(package_Anon_24_io_x_ppn),
    .io_x_u(package_Anon_24_io_x_u),
    .io_x_ae(package_Anon_24_io_x_ae),
    .io_x_sw(package_Anon_24_io_x_sw),
    .io_x_sx(package_Anon_24_io_x_sx),
    .io_x_sr(package_Anon_24_io_x_sr),
    .io_x_pw(package_Anon_24_io_x_pw),
    .io_x_px(package_Anon_24_io_x_px),
    .io_x_pr(package_Anon_24_io_x_pr),
    .io_x_pal(package_Anon_24_io_x_pal),
    .io_x_paa(package_Anon_24_io_x_paa),
    .io_x_eff(package_Anon_24_io_x_eff),
    .io_x_c(package_Anon_24_io_x_c),
    .io_y_ppn(package_Anon_24_io_y_ppn),
    .io_y_u(package_Anon_24_io_y_u),
    .io_y_ae(package_Anon_24_io_y_ae),
    .io_y_sw(package_Anon_24_io_y_sw),
    .io_y_sx(package_Anon_24_io_y_sx),
    .io_y_sr(package_Anon_24_io_y_sr),
    .io_y_pw(package_Anon_24_io_y_pw),
    .io_y_px(package_Anon_24_io_y_px),
    .io_y_pr(package_Anon_24_io_y_pr),
    .io_y_pal(package_Anon_24_io_y_pal),
    .io_y_paa(package_Anon_24_io_y_paa),
    .io_y_eff(package_Anon_24_io_y_eff),
    .io_y_c(package_Anon_24_io_y_c)
  );
  package_Anon package_Anon_25 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223114.4]
    .io_x_ppn(package_Anon_25_io_x_ppn),
    .io_x_u(package_Anon_25_io_x_u),
    .io_x_ae(package_Anon_25_io_x_ae),
    .io_x_sw(package_Anon_25_io_x_sw),
    .io_x_sx(package_Anon_25_io_x_sx),
    .io_x_sr(package_Anon_25_io_x_sr),
    .io_x_pw(package_Anon_25_io_x_pw),
    .io_x_px(package_Anon_25_io_x_px),
    .io_x_pr(package_Anon_25_io_x_pr),
    .io_x_pal(package_Anon_25_io_x_pal),
    .io_x_paa(package_Anon_25_io_x_paa),
    .io_x_eff(package_Anon_25_io_x_eff),
    .io_x_c(package_Anon_25_io_x_c),
    .io_y_ppn(package_Anon_25_io_y_ppn),
    .io_y_u(package_Anon_25_io_y_u),
    .io_y_ae(package_Anon_25_io_y_ae),
    .io_y_sw(package_Anon_25_io_y_sw),
    .io_y_sx(package_Anon_25_io_y_sx),
    .io_y_sr(package_Anon_25_io_y_sr),
    .io_y_pw(package_Anon_25_io_y_pw),
    .io_y_px(package_Anon_25_io_y_px),
    .io_y_pr(package_Anon_25_io_y_pr),
    .io_y_pal(package_Anon_25_io_y_pal),
    .io_y_paa(package_Anon_25_io_y_paa),
    .io_y_eff(package_Anon_25_io_y_eff),
    .io_y_c(package_Anon_25_io_y_c)
  );
  package_Anon package_Anon_26 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223154.4]
    .io_x_ppn(package_Anon_26_io_x_ppn),
    .io_x_u(package_Anon_26_io_x_u),
    .io_x_ae(package_Anon_26_io_x_ae),
    .io_x_sw(package_Anon_26_io_x_sw),
    .io_x_sx(package_Anon_26_io_x_sx),
    .io_x_sr(package_Anon_26_io_x_sr),
    .io_x_pw(package_Anon_26_io_x_pw),
    .io_x_px(package_Anon_26_io_x_px),
    .io_x_pr(package_Anon_26_io_x_pr),
    .io_x_pal(package_Anon_26_io_x_pal),
    .io_x_paa(package_Anon_26_io_x_paa),
    .io_x_eff(package_Anon_26_io_x_eff),
    .io_x_c(package_Anon_26_io_x_c),
    .io_y_ppn(package_Anon_26_io_y_ppn),
    .io_y_u(package_Anon_26_io_y_u),
    .io_y_ae(package_Anon_26_io_y_ae),
    .io_y_sw(package_Anon_26_io_y_sw),
    .io_y_sx(package_Anon_26_io_y_sx),
    .io_y_sr(package_Anon_26_io_y_sr),
    .io_y_pw(package_Anon_26_io_y_pw),
    .io_y_px(package_Anon_26_io_y_px),
    .io_y_pr(package_Anon_26_io_y_pr),
    .io_y_pal(package_Anon_26_io_y_pal),
    .io_y_paa(package_Anon_26_io_y_paa),
    .io_y_eff(package_Anon_26_io_y_eff),
    .io_y_c(package_Anon_26_io_y_c)
  );
  package_Anon package_Anon_27 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223195.4]
    .io_x_ppn(package_Anon_27_io_x_ppn),
    .io_x_u(package_Anon_27_io_x_u),
    .io_x_ae(package_Anon_27_io_x_ae),
    .io_x_sw(package_Anon_27_io_x_sw),
    .io_x_sx(package_Anon_27_io_x_sx),
    .io_x_sr(package_Anon_27_io_x_sr),
    .io_x_pw(package_Anon_27_io_x_pw),
    .io_x_px(package_Anon_27_io_x_px),
    .io_x_pr(package_Anon_27_io_x_pr),
    .io_x_pal(package_Anon_27_io_x_pal),
    .io_x_paa(package_Anon_27_io_x_paa),
    .io_x_eff(package_Anon_27_io_x_eff),
    .io_x_c(package_Anon_27_io_x_c),
    .io_y_ppn(package_Anon_27_io_y_ppn),
    .io_y_u(package_Anon_27_io_y_u),
    .io_y_ae(package_Anon_27_io_y_ae),
    .io_y_sw(package_Anon_27_io_y_sw),
    .io_y_sx(package_Anon_27_io_y_sx),
    .io_y_sr(package_Anon_27_io_y_sr),
    .io_y_pw(package_Anon_27_io_y_pw),
    .io_y_px(package_Anon_27_io_y_px),
    .io_y_pr(package_Anon_27_io_y_pr),
    .io_y_pal(package_Anon_27_io_y_pal),
    .io_y_paa(package_Anon_27_io_y_paa),
    .io_y_eff(package_Anon_27_io_y_eff),
    .io_y_c(package_Anon_27_io_y_c)
  );
  package_Anon package_Anon_28 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223236.4]
    .io_x_ppn(package_Anon_28_io_x_ppn),
    .io_x_u(package_Anon_28_io_x_u),
    .io_x_ae(package_Anon_28_io_x_ae),
    .io_x_sw(package_Anon_28_io_x_sw),
    .io_x_sx(package_Anon_28_io_x_sx),
    .io_x_sr(package_Anon_28_io_x_sr),
    .io_x_pw(package_Anon_28_io_x_pw),
    .io_x_px(package_Anon_28_io_x_px),
    .io_x_pr(package_Anon_28_io_x_pr),
    .io_x_pal(package_Anon_28_io_x_pal),
    .io_x_paa(package_Anon_28_io_x_paa),
    .io_x_eff(package_Anon_28_io_x_eff),
    .io_x_c(package_Anon_28_io_x_c),
    .io_y_ppn(package_Anon_28_io_y_ppn),
    .io_y_u(package_Anon_28_io_y_u),
    .io_y_ae(package_Anon_28_io_y_ae),
    .io_y_sw(package_Anon_28_io_y_sw),
    .io_y_sx(package_Anon_28_io_y_sx),
    .io_y_sr(package_Anon_28_io_y_sr),
    .io_y_pw(package_Anon_28_io_y_pw),
    .io_y_px(package_Anon_28_io_y_px),
    .io_y_pr(package_Anon_28_io_y_pr),
    .io_y_pal(package_Anon_28_io_y_pal),
    .io_y_paa(package_Anon_28_io_y_paa),
    .io_y_eff(package_Anon_28_io_y_eff),
    .io_y_c(package_Anon_28_io_y_c)
  );
  package_Anon package_Anon_29 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223277.4]
    .io_x_ppn(package_Anon_29_io_x_ppn),
    .io_x_u(package_Anon_29_io_x_u),
    .io_x_ae(package_Anon_29_io_x_ae),
    .io_x_sw(package_Anon_29_io_x_sw),
    .io_x_sx(package_Anon_29_io_x_sx),
    .io_x_sr(package_Anon_29_io_x_sr),
    .io_x_pw(package_Anon_29_io_x_pw),
    .io_x_px(package_Anon_29_io_x_px),
    .io_x_pr(package_Anon_29_io_x_pr),
    .io_x_pal(package_Anon_29_io_x_pal),
    .io_x_paa(package_Anon_29_io_x_paa),
    .io_x_eff(package_Anon_29_io_x_eff),
    .io_x_c(package_Anon_29_io_x_c),
    .io_y_ppn(package_Anon_29_io_y_ppn),
    .io_y_u(package_Anon_29_io_y_u),
    .io_y_ae(package_Anon_29_io_y_ae),
    .io_y_sw(package_Anon_29_io_y_sw),
    .io_y_sx(package_Anon_29_io_y_sx),
    .io_y_sr(package_Anon_29_io_y_sr),
    .io_y_pw(package_Anon_29_io_y_pw),
    .io_y_px(package_Anon_29_io_y_px),
    .io_y_pr(package_Anon_29_io_y_pr),
    .io_y_pal(package_Anon_29_io_y_pal),
    .io_y_paa(package_Anon_29_io_y_paa),
    .io_y_eff(package_Anon_29_io_y_eff),
    .io_y_c(package_Anon_29_io_y_c)
  );
  package_Anon package_Anon_30 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223318.4]
    .io_x_ppn(package_Anon_30_io_x_ppn),
    .io_x_u(package_Anon_30_io_x_u),
    .io_x_ae(package_Anon_30_io_x_ae),
    .io_x_sw(package_Anon_30_io_x_sw),
    .io_x_sx(package_Anon_30_io_x_sx),
    .io_x_sr(package_Anon_30_io_x_sr),
    .io_x_pw(package_Anon_30_io_x_pw),
    .io_x_px(package_Anon_30_io_x_px),
    .io_x_pr(package_Anon_30_io_x_pr),
    .io_x_pal(package_Anon_30_io_x_pal),
    .io_x_paa(package_Anon_30_io_x_paa),
    .io_x_eff(package_Anon_30_io_x_eff),
    .io_x_c(package_Anon_30_io_x_c),
    .io_y_ppn(package_Anon_30_io_y_ppn),
    .io_y_u(package_Anon_30_io_y_u),
    .io_y_ae(package_Anon_30_io_y_ae),
    .io_y_sw(package_Anon_30_io_y_sw),
    .io_y_sx(package_Anon_30_io_y_sx),
    .io_y_sr(package_Anon_30_io_y_sr),
    .io_y_pw(package_Anon_30_io_y_pw),
    .io_y_px(package_Anon_30_io_y_px),
    .io_y_pr(package_Anon_30_io_y_pr),
    .io_y_pal(package_Anon_30_io_y_pal),
    .io_y_paa(package_Anon_30_io_y_paa),
    .io_y_eff(package_Anon_30_io_y_eff),
    .io_y_c(package_Anon_30_io_y_c)
  );
  package_Anon package_Anon_31 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223359.4]
    .io_x_ppn(package_Anon_31_io_x_ppn),
    .io_x_u(package_Anon_31_io_x_u),
    .io_x_ae(package_Anon_31_io_x_ae),
    .io_x_sw(package_Anon_31_io_x_sw),
    .io_x_sx(package_Anon_31_io_x_sx),
    .io_x_sr(package_Anon_31_io_x_sr),
    .io_x_pw(package_Anon_31_io_x_pw),
    .io_x_px(package_Anon_31_io_x_px),
    .io_x_pr(package_Anon_31_io_x_pr),
    .io_x_pal(package_Anon_31_io_x_pal),
    .io_x_paa(package_Anon_31_io_x_paa),
    .io_x_eff(package_Anon_31_io_x_eff),
    .io_x_c(package_Anon_31_io_x_c),
    .io_y_ppn(package_Anon_31_io_y_ppn),
    .io_y_u(package_Anon_31_io_y_u),
    .io_y_ae(package_Anon_31_io_y_ae),
    .io_y_sw(package_Anon_31_io_y_sw),
    .io_y_sx(package_Anon_31_io_y_sx),
    .io_y_sr(package_Anon_31_io_y_sr),
    .io_y_pw(package_Anon_31_io_y_pw),
    .io_y_px(package_Anon_31_io_y_px),
    .io_y_pr(package_Anon_31_io_y_pr),
    .io_y_pal(package_Anon_31_io_y_pal),
    .io_y_paa(package_Anon_31_io_y_paa),
    .io_y_eff(package_Anon_31_io_y_eff),
    .io_y_c(package_Anon_31_io_y_c)
  );
  package_Anon package_Anon_32 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223400.4]
    .io_x_ppn(package_Anon_32_io_x_ppn),
    .io_x_u(package_Anon_32_io_x_u),
    .io_x_ae(package_Anon_32_io_x_ae),
    .io_x_sw(package_Anon_32_io_x_sw),
    .io_x_sx(package_Anon_32_io_x_sx),
    .io_x_sr(package_Anon_32_io_x_sr),
    .io_x_pw(package_Anon_32_io_x_pw),
    .io_x_px(package_Anon_32_io_x_px),
    .io_x_pr(package_Anon_32_io_x_pr),
    .io_x_pal(package_Anon_32_io_x_pal),
    .io_x_paa(package_Anon_32_io_x_paa),
    .io_x_eff(package_Anon_32_io_x_eff),
    .io_x_c(package_Anon_32_io_x_c),
    .io_y_ppn(package_Anon_32_io_y_ppn),
    .io_y_u(package_Anon_32_io_y_u),
    .io_y_ae(package_Anon_32_io_y_ae),
    .io_y_sw(package_Anon_32_io_y_sw),
    .io_y_sx(package_Anon_32_io_y_sx),
    .io_y_sr(package_Anon_32_io_y_sr),
    .io_y_pw(package_Anon_32_io_y_pw),
    .io_y_px(package_Anon_32_io_y_px),
    .io_y_pr(package_Anon_32_io_y_pr),
    .io_y_pal(package_Anon_32_io_y_pal),
    .io_y_paa(package_Anon_32_io_y_paa),
    .io_y_eff(package_Anon_32_io_y_eff),
    .io_y_c(package_Anon_32_io_y_c)
  );
  package_Anon package_Anon_33 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223441.4]
    .io_x_ppn(package_Anon_33_io_x_ppn),
    .io_x_u(package_Anon_33_io_x_u),
    .io_x_ae(package_Anon_33_io_x_ae),
    .io_x_sw(package_Anon_33_io_x_sw),
    .io_x_sx(package_Anon_33_io_x_sx),
    .io_x_sr(package_Anon_33_io_x_sr),
    .io_x_pw(package_Anon_33_io_x_pw),
    .io_x_px(package_Anon_33_io_x_px),
    .io_x_pr(package_Anon_33_io_x_pr),
    .io_x_pal(package_Anon_33_io_x_pal),
    .io_x_paa(package_Anon_33_io_x_paa),
    .io_x_eff(package_Anon_33_io_x_eff),
    .io_x_c(package_Anon_33_io_x_c),
    .io_y_ppn(package_Anon_33_io_y_ppn),
    .io_y_u(package_Anon_33_io_y_u),
    .io_y_ae(package_Anon_33_io_y_ae),
    .io_y_sw(package_Anon_33_io_y_sw),
    .io_y_sx(package_Anon_33_io_y_sx),
    .io_y_sr(package_Anon_33_io_y_sr),
    .io_y_pw(package_Anon_33_io_y_pw),
    .io_y_px(package_Anon_33_io_y_px),
    .io_y_pr(package_Anon_33_io_y_pr),
    .io_y_pal(package_Anon_33_io_y_pal),
    .io_y_paa(package_Anon_33_io_y_paa),
    .io_y_eff(package_Anon_33_io_y_eff),
    .io_y_c(package_Anon_33_io_y_c)
  );
  package_Anon package_Anon_34 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223482.4]
    .io_x_ppn(package_Anon_34_io_x_ppn),
    .io_x_u(package_Anon_34_io_x_u),
    .io_x_ae(package_Anon_34_io_x_ae),
    .io_x_sw(package_Anon_34_io_x_sw),
    .io_x_sx(package_Anon_34_io_x_sx),
    .io_x_sr(package_Anon_34_io_x_sr),
    .io_x_pw(package_Anon_34_io_x_pw),
    .io_x_px(package_Anon_34_io_x_px),
    .io_x_pr(package_Anon_34_io_x_pr),
    .io_x_pal(package_Anon_34_io_x_pal),
    .io_x_paa(package_Anon_34_io_x_paa),
    .io_x_eff(package_Anon_34_io_x_eff),
    .io_x_c(package_Anon_34_io_x_c),
    .io_y_ppn(package_Anon_34_io_y_ppn),
    .io_y_u(package_Anon_34_io_y_u),
    .io_y_ae(package_Anon_34_io_y_ae),
    .io_y_sw(package_Anon_34_io_y_sw),
    .io_y_sx(package_Anon_34_io_y_sx),
    .io_y_sr(package_Anon_34_io_y_sr),
    .io_y_pw(package_Anon_34_io_y_pw),
    .io_y_px(package_Anon_34_io_y_px),
    .io_y_pr(package_Anon_34_io_y_pr),
    .io_y_pal(package_Anon_34_io_y_pal),
    .io_y_paa(package_Anon_34_io_y_paa),
    .io_y_eff(package_Anon_34_io_y_eff),
    .io_y_c(package_Anon_34_io_y_c)
  );
  package_Anon package_Anon_35 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223522.4]
    .io_x_ppn(package_Anon_35_io_x_ppn),
    .io_x_u(package_Anon_35_io_x_u),
    .io_x_ae(package_Anon_35_io_x_ae),
    .io_x_sw(package_Anon_35_io_x_sw),
    .io_x_sx(package_Anon_35_io_x_sx),
    .io_x_sr(package_Anon_35_io_x_sr),
    .io_x_pw(package_Anon_35_io_x_pw),
    .io_x_px(package_Anon_35_io_x_px),
    .io_x_pr(package_Anon_35_io_x_pr),
    .io_x_pal(package_Anon_35_io_x_pal),
    .io_x_paa(package_Anon_35_io_x_paa),
    .io_x_eff(package_Anon_35_io_x_eff),
    .io_x_c(package_Anon_35_io_x_c),
    .io_y_ppn(package_Anon_35_io_y_ppn),
    .io_y_u(package_Anon_35_io_y_u),
    .io_y_ae(package_Anon_35_io_y_ae),
    .io_y_sw(package_Anon_35_io_y_sw),
    .io_y_sx(package_Anon_35_io_y_sx),
    .io_y_sr(package_Anon_35_io_y_sr),
    .io_y_pw(package_Anon_35_io_y_pw),
    .io_y_px(package_Anon_35_io_y_px),
    .io_y_pr(package_Anon_35_io_y_pr),
    .io_y_pal(package_Anon_35_io_y_pal),
    .io_y_paa(package_Anon_35_io_y_paa),
    .io_y_eff(package_Anon_35_io_y_eff),
    .io_y_c(package_Anon_35_io_y_c)
  );
  package_Anon package_Anon_36 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223562.4]
    .io_x_ppn(package_Anon_36_io_x_ppn),
    .io_x_u(package_Anon_36_io_x_u),
    .io_x_ae(package_Anon_36_io_x_ae),
    .io_x_sw(package_Anon_36_io_x_sw),
    .io_x_sx(package_Anon_36_io_x_sx),
    .io_x_sr(package_Anon_36_io_x_sr),
    .io_x_pw(package_Anon_36_io_x_pw),
    .io_x_px(package_Anon_36_io_x_px),
    .io_x_pr(package_Anon_36_io_x_pr),
    .io_x_pal(package_Anon_36_io_x_pal),
    .io_x_paa(package_Anon_36_io_x_paa),
    .io_x_eff(package_Anon_36_io_x_eff),
    .io_x_c(package_Anon_36_io_x_c),
    .io_y_ppn(package_Anon_36_io_y_ppn),
    .io_y_u(package_Anon_36_io_y_u),
    .io_y_ae(package_Anon_36_io_y_ae),
    .io_y_sw(package_Anon_36_io_y_sw),
    .io_y_sx(package_Anon_36_io_y_sx),
    .io_y_sr(package_Anon_36_io_y_sr),
    .io_y_pw(package_Anon_36_io_y_pw),
    .io_y_px(package_Anon_36_io_y_px),
    .io_y_pr(package_Anon_36_io_y_pr),
    .io_y_pal(package_Anon_36_io_y_pal),
    .io_y_paa(package_Anon_36_io_y_paa),
    .io_y_eff(package_Anon_36_io_y_eff),
    .io_y_c(package_Anon_36_io_y_c)
  );
  package_Anon package_Anon_37 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223602.4]
    .io_x_ppn(package_Anon_37_io_x_ppn),
    .io_x_u(package_Anon_37_io_x_u),
    .io_x_ae(package_Anon_37_io_x_ae),
    .io_x_sw(package_Anon_37_io_x_sw),
    .io_x_sx(package_Anon_37_io_x_sx),
    .io_x_sr(package_Anon_37_io_x_sr),
    .io_x_pw(package_Anon_37_io_x_pw),
    .io_x_px(package_Anon_37_io_x_px),
    .io_x_pr(package_Anon_37_io_x_pr),
    .io_x_pal(package_Anon_37_io_x_pal),
    .io_x_paa(package_Anon_37_io_x_paa),
    .io_x_eff(package_Anon_37_io_x_eff),
    .io_x_c(package_Anon_37_io_x_c),
    .io_y_ppn(package_Anon_37_io_y_ppn),
    .io_y_u(package_Anon_37_io_y_u),
    .io_y_ae(package_Anon_37_io_y_ae),
    .io_y_sw(package_Anon_37_io_y_sw),
    .io_y_sx(package_Anon_37_io_y_sx),
    .io_y_sr(package_Anon_37_io_y_sr),
    .io_y_pw(package_Anon_37_io_y_pw),
    .io_y_px(package_Anon_37_io_y_px),
    .io_y_pr(package_Anon_37_io_y_pr),
    .io_y_pal(package_Anon_37_io_y_pal),
    .io_y_paa(package_Anon_37_io_y_paa),
    .io_y_eff(package_Anon_37_io_y_eff),
    .io_y_c(package_Anon_37_io_y_c)
  );
  package_Anon package_Anon_38 ( // @[package.scala 213:21:chipyard.TestHarness.RocketConfig.fir@223642.4]
    .io_x_ppn(package_Anon_38_io_x_ppn),
    .io_x_u(package_Anon_38_io_x_u),
    .io_x_ae(package_Anon_38_io_x_ae),
    .io_x_sw(package_Anon_38_io_x_sw),
    .io_x_sx(package_Anon_38_io_x_sx),
    .io_x_sr(package_Anon_38_io_x_sr),
    .io_x_pw(package_Anon_38_io_x_pw),
    .io_x_px(package_Anon_38_io_x_px),
    .io_x_pr(package_Anon_38_io_x_pr),
    .io_x_pal(package_Anon_38_io_x_pal),
    .io_x_paa(package_Anon_38_io_x_paa),
    .io_x_eff(package_Anon_38_io_x_eff),
    .io_x_c(package_Anon_38_io_x_c),
    .io_y_ppn(package_Anon_38_io_y_ppn),
    .io_y_u(package_Anon_38_io_y_u),
    .io_y_ae(package_Anon_38_io_y_ae),
    .io_y_sw(package_Anon_38_io_y_sw),
    .io_y_sx(package_Anon_38_io_y_sx),
    .io_y_sr(package_Anon_38_io_y_sr),
    .io_y_pw(package_Anon_38_io_y_pw),
    .io_y_px(package_Anon_38_io_y_px),
    .io_y_pr(package_Anon_38_io_y_pr),
    .io_y_pal(package_Anon_38_io_y_pal),
    .io_y_paa(package_Anon_38_io_y_paa),
    .io_y_eff(package_Anon_38_io_y_eff),
    .io_y_c(package_Anon_38_io_y_c)
  );
  assign priv_s = io_ptw_status_prv[0]; // @[TLB.scala 176:20:chipyard.TestHarness.RocketConfig.fir@220847.4]
  assign priv_uses_vm = io_ptw_status_prv <= 2'h1; // @[TLB.scala 177:27:chipyard.TestHarness.RocketConfig.fir@220848.4]
  assign vm_enabled = io_ptw_ptbr_mode[3] & priv_uses_vm; // @[TLB.scala 178:83:chipyard.TestHarness.RocketConfig.fir@220851.4]
  assign vpn = io_req_bits_vaddr[38:12]; // @[TLB.scala 181:30:chipyard.TestHarness.RocketConfig.fir@220854.4]
  assign refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[TLB.scala 182:44:chipyard.TestHarness.RocketConfig.fir@220855.4]
  assign _T_4 = state == 2'h1; // @[package.scala 15:47:chipyard.TestHarness.RocketConfig.fir@220857.4]
  assign _T_5 = state == 2'h3; // @[package.scala 15:47:chipyard.TestHarness.RocketConfig.fir@220858.4]
  assign invalidate_refill = _T_4 | _T_5; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@220859.4]
  assign _T_25 = special_entry_level < 2'h1; // @[TLB.scala 107:28:chipyard.TestHarness.RocketConfig.fir@220902.4]
  assign _T_27 = _T_25 ? vpn : 27'h0; // @[TLB.scala 108:28:chipyard.TestHarness.RocketConfig.fir@220904.4]
  assign _GEN_950 = {{7'd0}, package_Anon_io_y_ppn}; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@220905.4]
  assign _T_28 = _T_27 | _GEN_950; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@220905.4]
  assign _T_31 = special_entry_level < 2'h2; // @[TLB.scala 107:28:chipyard.TestHarness.RocketConfig.fir@220908.4]
  assign _T_33 = _T_31 ? vpn : 27'h0; // @[TLB.scala 108:28:chipyard.TestHarness.RocketConfig.fir@220910.4]
  assign _T_34 = _T_33 | _GEN_950; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@220911.4]
  assign _T_36 = {package_Anon_io_y_ppn[19:18],_T_28[17:9],_T_34[8:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@220913.4]
  assign _T_38 = vm_enabled ? {{8'd0}, _T_36} : io_req_bits_vaddr[39:12]; // @[TLB.scala 186:20:chipyard.TestHarness.RocketConfig.fir@220915.4]
  assign mpu_ppn = io_ptw_resp_valid ? {{8'd0}, refill_ppn} : _T_38; // @[TLB.scala 185:20:chipyard.TestHarness.RocketConfig.fir@220916.4]
  assign mpu_physaddr = {mpu_ppn,io_req_bits_vaddr[11:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@220918.4]
  assign _T_42 = {io_ptw_status_debug,io_ptw_status_prv}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@220921.4]
  assign mpu_priv = io_ptw_resp_valid ? 3'h1 : _T_42; // @[TLB.scala 188:27:chipyard.TestHarness.RocketConfig.fir@220922.4]
  assign _T_43 = mpu_physaddr ^ 40'h3000; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220938.4]
  assign _T_44 = {1'b0,$signed(_T_43)}; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220939.4]
  assign _T_46 = $signed(_T_44) & -41'sh1000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220941.4]
  assign _T_47 = $signed(_T_46) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220942.4]
  assign _T_48 = mpu_physaddr ^ 40'h2010000; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220943.4]
  assign _T_49 = {1'b0,$signed(_T_48)}; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220944.4]
  assign _T_51 = $signed(_T_49) & -41'sh1000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220946.4]
  assign _T_52 = $signed(_T_51) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220947.4]
  assign _T_53 = mpu_physaddr ^ 40'h54000000; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220948.4]
  assign _T_54 = {1'b0,$signed(_T_53)}; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220949.4]
  assign _T_56 = $signed(_T_54) & -41'sh1000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220951.4]
  assign _T_57 = $signed(_T_56) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220952.4]
  assign _T_58 = mpu_physaddr ^ 40'hc000000; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220953.4]
  assign _T_59 = {1'b0,$signed(_T_58)}; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220954.4]
  assign _T_61 = $signed(_T_59) & -41'sh4000000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220956.4]
  assign _T_62 = $signed(_T_61) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220957.4]
  assign _T_63 = mpu_physaddr ^ 40'h2000000; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220958.4]
  assign _T_64 = {1'b0,$signed(_T_63)}; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220959.4]
  assign _T_66 = $signed(_T_64) & -41'sh10000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220961.4]
  assign _T_67 = $signed(_T_66) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220962.4]
  assign _T_69 = {1'b0,$signed(mpu_physaddr)}; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220964.4]
  assign _T_71 = $signed(_T_69) & -41'sh1000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220966.4]
  assign _T_72 = $signed(_T_71) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220967.4]
  assign _T_73 = mpu_physaddr ^ 40'h10000; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220968.4]
  assign _T_74 = {1'b0,$signed(_T_73)}; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220969.4]
  assign _T_76 = $signed(_T_74) & -41'sh10000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220971.4]
  assign _T_77 = $signed(_T_76) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220972.4]
  assign _T_78 = mpu_physaddr ^ 40'h80000000; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@220973.4]
  assign _T_79 = {1'b0,$signed(_T_78)}; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@220974.4]
  assign _T_81 = $signed(_T_79) & -41'sh10000000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@220976.4]
  assign _T_82 = $signed(_T_81) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@220977.4]
  assign _T_84 = _T_47 | _T_52; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220988.4]
  assign _T_85 = _T_84 | _T_57; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220989.4]
  assign _T_86 = _T_85 | _T_62; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220990.4]
  assign _T_87 = _T_86 | _T_67; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220991.4]
  assign _T_88 = _T_87 | _T_72; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220992.4]
  assign _T_89 = _T_88 | _T_77; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220993.4]
  assign legal_address = _T_89 | _T_82; // @[TLB.scala 194:67:chipyard.TestHarness.RocketConfig.fir@220994.4]
  assign _T_98 = $signed(_T_79) & 41'sh80000000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221003.4]
  assign _T_99 = $signed(_T_98) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221004.4]
  assign cacheable = legal_address & _T_99; // @[TLB.scala 196:19:chipyard.TestHarness.RocketConfig.fir@221010.4]
  assign _T_163 = $signed(_T_69) & 41'sh86000000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221071.4]
  assign _T_164 = $signed(_T_163) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221072.4]
  assign _T_171 = _T_164 | _T_99; // @[TLBPermissions.scala 82:66:chipyard.TestHarness.RocketConfig.fir@221079.4]
  assign _T_192 = mpu_priv <= 3'h3; // @[TLB.scala 199:39:chipyard.TestHarness.RocketConfig.fir@221100.4]
  assign deny_access_to_debug = _T_192 & _T_72; // @[TLB.scala 199:48:chipyard.TestHarness.RocketConfig.fir@221106.4]
  assign _T_204 = ~deny_access_to_debug; // @[TLB.scala 200:44:chipyard.TestHarness.RocketConfig.fir@221113.4]
  assign _T_205 = legal_address & _T_204; // @[TLB.scala 200:41:chipyard.TestHarness.RocketConfig.fir@221114.4]
  assign prot_r = _T_205 & pmp_io_r; // @[TLB.scala 200:66:chipyard.TestHarness.RocketConfig.fir@221115.4]
  assign _T_209 = $signed(_T_69) & 41'sh82010000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221119.4]
  assign _T_210 = $signed(_T_209) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221120.4]
  assign _T_214 = $signed(_T_64) & 41'sh86000000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221124.4]
  assign _T_215 = $signed(_T_214) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221125.4]
  assign _T_216 = mpu_physaddr ^ 40'h4000000; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@221126.4]
  assign _T_217 = {1'b0,$signed(_T_216)}; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@221127.4]
  assign _T_219 = $signed(_T_217) & 41'sh84000000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221129.4]
  assign _T_220 = $signed(_T_219) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221130.4]
  assign _T_226 = _T_210 | _T_215; // @[Parameters.scala 528:89:chipyard.TestHarness.RocketConfig.fir@221136.4]
  assign _T_227 = _T_226 | _T_220; // @[Parameters.scala 528:89:chipyard.TestHarness.RocketConfig.fir@221137.4]
  assign _T_228 = _T_227 | _T_99; // @[Parameters.scala 528:89:chipyard.TestHarness.RocketConfig.fir@221138.4]
  assign _T_238 = legal_address & _T_228; // @[TLB.scala 196:19:chipyard.TestHarness.RocketConfig.fir@221149.4]
  assign _T_240 = _T_238 & _T_204; // @[TLB.scala 201:45:chipyard.TestHarness.RocketConfig.fir@221151.4]
  assign prot_w = _T_240 & pmp_io_w; // @[TLB.scala 201:70:chipyard.TestHarness.RocketConfig.fir@221152.4]
  assign _T_337 = legal_address & _T_171; // @[TLB.scala 196:19:chipyard.TestHarness.RocketConfig.fir@221254.4]
  assign _T_339 = _T_337 & _T_204; // @[TLB.scala 204:40:chipyard.TestHarness.RocketConfig.fir@221256.4]
  assign prot_x = _T_339 & pmp_io_x; // @[TLB.scala 204:65:chipyard.TestHarness.RocketConfig.fir@221257.4]
  assign _T_360 = $signed(_T_49) & 41'sh86012000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221278.4]
  assign _T_361 = $signed(_T_360) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221279.4]
  assign _T_365 = $signed(_T_69) & 41'sh82012000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221283.4]
  assign _T_366 = $signed(_T_365) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221284.4]
  assign _T_375 = $signed(_T_64) & 41'sh86010000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@221293.4]
  assign _T_376 = $signed(_T_375) == 41'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@221294.4]
  assign _T_377 = _T_361 | _T_366; // @[Parameters.scala 528:89:chipyard.TestHarness.RocketConfig.fir@221295.4]
  assign _T_378 = _T_377 | _T_220; // @[Parameters.scala 528:89:chipyard.TestHarness.RocketConfig.fir@221296.4]
  assign _T_379 = _T_378 | _T_376; // @[Parameters.scala 528:89:chipyard.TestHarness.RocketConfig.fir@221297.4]
  assign prot_eff = legal_address & _T_379; // @[TLB.scala 196:19:chipyard.TestHarness.RocketConfig.fir@221303.4]
  assign _T_384 = sectored_entries_0_valid_0 | sectored_entries_0_valid_1; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221304.4]
  assign _T_385 = _T_384 | sectored_entries_0_valid_2; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221305.4]
  assign _T_386 = _T_385 | sectored_entries_0_valid_3; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221306.4]
  assign _T_387 = sectored_entries_0_tag ^ vpn; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221307.4]
  assign _T_389 = _T_387[26:2] == 25'h0; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221309.4]
  assign sector_hits_0 = _T_386 & _T_389; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221310.4]
  assign _T_390 = sectored_entries_1_valid_0 | sectored_entries_1_valid_1; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221311.4]
  assign _T_391 = _T_390 | sectored_entries_1_valid_2; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221312.4]
  assign _T_392 = _T_391 | sectored_entries_1_valid_3; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221313.4]
  assign _T_393 = sectored_entries_1_tag ^ vpn; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221314.4]
  assign _T_395 = _T_393[26:2] == 25'h0; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221316.4]
  assign sector_hits_1 = _T_392 & _T_395; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221317.4]
  assign _T_396 = sectored_entries_2_valid_0 | sectored_entries_2_valid_1; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221318.4]
  assign _T_397 = _T_396 | sectored_entries_2_valid_2; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221319.4]
  assign _T_398 = _T_397 | sectored_entries_2_valid_3; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221320.4]
  assign _T_399 = sectored_entries_2_tag ^ vpn; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221321.4]
  assign _T_401 = _T_399[26:2] == 25'h0; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221323.4]
  assign sector_hits_2 = _T_398 & _T_401; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221324.4]
  assign _T_402 = sectored_entries_3_valid_0 | sectored_entries_3_valid_1; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221325.4]
  assign _T_403 = _T_402 | sectored_entries_3_valid_2; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221326.4]
  assign _T_404 = _T_403 | sectored_entries_3_valid_3; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221327.4]
  assign _T_405 = sectored_entries_3_tag ^ vpn; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221328.4]
  assign _T_407 = _T_405[26:2] == 25'h0; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221330.4]
  assign sector_hits_3 = _T_404 & _T_407; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221331.4]
  assign _T_408 = sectored_entries_4_valid_0 | sectored_entries_4_valid_1; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221332.4]
  assign _T_409 = _T_408 | sectored_entries_4_valid_2; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221333.4]
  assign _T_410 = _T_409 | sectored_entries_4_valid_3; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221334.4]
  assign _T_411 = sectored_entries_4_tag ^ vpn; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221335.4]
  assign _T_413 = _T_411[26:2] == 25'h0; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221337.4]
  assign sector_hits_4 = _T_410 & _T_413; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221338.4]
  assign _T_414 = sectored_entries_5_valid_0 | sectored_entries_5_valid_1; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221339.4]
  assign _T_415 = _T_414 | sectored_entries_5_valid_2; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221340.4]
  assign _T_416 = _T_415 | sectored_entries_5_valid_3; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221341.4]
  assign _T_417 = sectored_entries_5_tag ^ vpn; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221342.4]
  assign _T_419 = _T_417[26:2] == 25'h0; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221344.4]
  assign sector_hits_5 = _T_416 & _T_419; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221345.4]
  assign _T_420 = sectored_entries_6_valid_0 | sectored_entries_6_valid_1; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221346.4]
  assign _T_421 = _T_420 | sectored_entries_6_valid_2; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221347.4]
  assign _T_422 = _T_421 | sectored_entries_6_valid_3; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221348.4]
  assign _T_423 = sectored_entries_6_tag ^ vpn; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221349.4]
  assign _T_425 = _T_423[26:2] == 25'h0; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221351.4]
  assign sector_hits_6 = _T_422 & _T_425; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221352.4]
  assign _T_426 = sectored_entries_7_valid_0 | sectored_entries_7_valid_1; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221353.4]
  assign _T_427 = _T_426 | sectored_entries_7_valid_2; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221354.4]
  assign _T_428 = _T_427 | sectored_entries_7_valid_3; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@221355.4]
  assign _T_429 = sectored_entries_7_tag ^ vpn; // @[TLB.scala 87:41:chipyard.TestHarness.RocketConfig.fir@221356.4]
  assign _T_431 = _T_429[26:2] == 25'h0; // @[TLB.scala 87:66:chipyard.TestHarness.RocketConfig.fir@221358.4]
  assign sector_hits_7 = _T_428 & _T_431; // @[TLB.scala 86:40:chipyard.TestHarness.RocketConfig.fir@221359.4]
  assign _T_436 = superpage_entries_0_tag[26:18] == vpn[26:18]; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221364.4]
  assign _T_438 = superpage_entries_0_valid_0 & _T_436; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221366.4]
  assign _T_439 = superpage_entries_0_level < 2'h1; // @[TLB.scala 93:28:chipyard.TestHarness.RocketConfig.fir@221367.4]
  assign _T_443 = superpage_entries_0_tag[17:9] == vpn[17:9]; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221371.4]
  assign _T_444 = _T_439 | _T_443; // @[TLB.scala 94:40:chipyard.TestHarness.RocketConfig.fir@221372.4]
  assign superpage_hits_0 = _T_438 & _T_444; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221373.4]
  assign _T_456 = superpage_entries_1_tag[26:18] == vpn[26:18]; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221385.4]
  assign _T_458 = superpage_entries_1_valid_0 & _T_456; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221387.4]
  assign _T_459 = superpage_entries_1_level < 2'h1; // @[TLB.scala 93:28:chipyard.TestHarness.RocketConfig.fir@221388.4]
  assign _T_463 = superpage_entries_1_tag[17:9] == vpn[17:9]; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221392.4]
  assign _T_464 = _T_459 | _T_463; // @[TLB.scala 94:40:chipyard.TestHarness.RocketConfig.fir@221393.4]
  assign superpage_hits_1 = _T_458 & _T_464; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221394.4]
  assign _T_476 = superpage_entries_2_tag[26:18] == vpn[26:18]; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221406.4]
  assign _T_478 = superpage_entries_2_valid_0 & _T_476; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221408.4]
  assign _T_479 = superpage_entries_2_level < 2'h1; // @[TLB.scala 93:28:chipyard.TestHarness.RocketConfig.fir@221409.4]
  assign _T_483 = superpage_entries_2_tag[17:9] == vpn[17:9]; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221413.4]
  assign _T_484 = _T_479 | _T_483; // @[TLB.scala 94:40:chipyard.TestHarness.RocketConfig.fir@221414.4]
  assign superpage_hits_2 = _T_478 & _T_484; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221415.4]
  assign _T_496 = superpage_entries_3_tag[26:18] == vpn[26:18]; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221427.4]
  assign _T_498 = superpage_entries_3_valid_0 & _T_496; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221429.4]
  assign _T_499 = superpage_entries_3_level < 2'h1; // @[TLB.scala 93:28:chipyard.TestHarness.RocketConfig.fir@221430.4]
  assign _T_503 = superpage_entries_3_tag[17:9] == vpn[17:9]; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221434.4]
  assign _T_504 = _T_499 | _T_503; // @[TLB.scala 94:40:chipyard.TestHarness.RocketConfig.fir@221435.4]
  assign superpage_hits_3 = _T_498 & _T_504; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221436.4]
  assign _GEN_1 = 2'h1 == vpn[1:0] ? sectored_entries_0_valid_1 : sectored_entries_0_valid_0; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221448.4]
  assign _GEN_2 = 2'h2 == vpn[1:0] ? sectored_entries_0_valid_2 : _GEN_1; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221448.4]
  assign _GEN_3 = 2'h3 == vpn[1:0] ? sectored_entries_0_valid_3 : _GEN_2; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221448.4]
  assign _T_516 = _GEN_3 & _T_389; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221448.4]
  assign hitsVec_0 = vm_enabled & _T_516; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221449.4]
  assign _GEN_5 = 2'h1 == vpn[1:0] ? sectored_entries_1_valid_1 : sectored_entries_1_valid_0; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221454.4]
  assign _GEN_6 = 2'h2 == vpn[1:0] ? sectored_entries_1_valid_2 : _GEN_5; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221454.4]
  assign _GEN_7 = 2'h3 == vpn[1:0] ? sectored_entries_1_valid_3 : _GEN_6; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221454.4]
  assign _T_521 = _GEN_7 & _T_395; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221454.4]
  assign hitsVec_1 = vm_enabled & _T_521; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221455.4]
  assign _GEN_9 = 2'h1 == vpn[1:0] ? sectored_entries_2_valid_1 : sectored_entries_2_valid_0; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221460.4]
  assign _GEN_10 = 2'h2 == vpn[1:0] ? sectored_entries_2_valid_2 : _GEN_9; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221460.4]
  assign _GEN_11 = 2'h3 == vpn[1:0] ? sectored_entries_2_valid_3 : _GEN_10; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221460.4]
  assign _T_526 = _GEN_11 & _T_401; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221460.4]
  assign hitsVec_2 = vm_enabled & _T_526; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221461.4]
  assign _GEN_13 = 2'h1 == vpn[1:0] ? sectored_entries_3_valid_1 : sectored_entries_3_valid_0; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221466.4]
  assign _GEN_14 = 2'h2 == vpn[1:0] ? sectored_entries_3_valid_2 : _GEN_13; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221466.4]
  assign _GEN_15 = 2'h3 == vpn[1:0] ? sectored_entries_3_valid_3 : _GEN_14; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221466.4]
  assign _T_531 = _GEN_15 & _T_407; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221466.4]
  assign hitsVec_3 = vm_enabled & _T_531; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221467.4]
  assign _GEN_17 = 2'h1 == vpn[1:0] ? sectored_entries_4_valid_1 : sectored_entries_4_valid_0; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221472.4]
  assign _GEN_18 = 2'h2 == vpn[1:0] ? sectored_entries_4_valid_2 : _GEN_17; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221472.4]
  assign _GEN_19 = 2'h3 == vpn[1:0] ? sectored_entries_4_valid_3 : _GEN_18; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221472.4]
  assign _T_536 = _GEN_19 & _T_413; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221472.4]
  assign hitsVec_4 = vm_enabled & _T_536; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221473.4]
  assign _GEN_21 = 2'h1 == vpn[1:0] ? sectored_entries_5_valid_1 : sectored_entries_5_valid_0; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221478.4]
  assign _GEN_22 = 2'h2 == vpn[1:0] ? sectored_entries_5_valid_2 : _GEN_21; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221478.4]
  assign _GEN_23 = 2'h3 == vpn[1:0] ? sectored_entries_5_valid_3 : _GEN_22; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221478.4]
  assign _T_541 = _GEN_23 & _T_419; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221478.4]
  assign hitsVec_5 = vm_enabled & _T_541; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221479.4]
  assign _GEN_25 = 2'h1 == vpn[1:0] ? sectored_entries_6_valid_1 : sectored_entries_6_valid_0; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221484.4]
  assign _GEN_26 = 2'h2 == vpn[1:0] ? sectored_entries_6_valid_2 : _GEN_25; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221484.4]
  assign _GEN_27 = 2'h3 == vpn[1:0] ? sectored_entries_6_valid_3 : _GEN_26; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221484.4]
  assign _T_546 = _GEN_27 & _T_425; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221484.4]
  assign hitsVec_6 = vm_enabled & _T_546; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221485.4]
  assign _GEN_29 = 2'h1 == vpn[1:0] ? sectored_entries_7_valid_1 : sectored_entries_7_valid_0; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221490.4]
  assign _GEN_30 = 2'h2 == vpn[1:0] ? sectored_entries_7_valid_2 : _GEN_29; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221490.4]
  assign _GEN_31 = 2'h3 == vpn[1:0] ? sectored_entries_7_valid_3 : _GEN_30; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221490.4]
  assign _T_551 = _GEN_31 & _T_431; // @[TLB.scala 99:18:chipyard.TestHarness.RocketConfig.fir@221490.4]
  assign hitsVec_7 = vm_enabled & _T_551; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221491.4]
  assign hitsVec_8 = vm_enabled & superpage_hits_0; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221513.4]
  assign hitsVec_9 = vm_enabled & superpage_hits_1; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221535.4]
  assign hitsVec_10 = vm_enabled & superpage_hits_2; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221557.4]
  assign hitsVec_11 = vm_enabled & superpage_hits_3; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221579.4]
  assign _T_640 = special_entry_tag[26:18] == vpn[26:18]; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221584.4]
  assign _T_642 = special_entry_valid_0 & _T_640; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221586.4]
  assign _T_647 = special_entry_tag[17:9] == vpn[17:9]; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221591.4]
  assign _T_648 = _T_25 | _T_647; // @[TLB.scala 94:40:chipyard.TestHarness.RocketConfig.fir@221592.4]
  assign _T_649 = _T_642 & _T_648; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221593.4]
  assign _T_654 = special_entry_tag[8:0] == vpn[8:0]; // @[TLB.scala 94:77:chipyard.TestHarness.RocketConfig.fir@221598.4]
  assign _T_655 = _T_31 | _T_654; // @[TLB.scala 94:40:chipyard.TestHarness.RocketConfig.fir@221599.4]
  assign _T_656 = _T_649 & _T_655; // @[TLB.scala 94:29:chipyard.TestHarness.RocketConfig.fir@221600.4]
  assign hitsVec_12 = vm_enabled & _T_656; // @[TLB.scala 209:44:chipyard.TestHarness.RocketConfig.fir@221601.4]
  assign _T_661 = {hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@221606.4]
  assign real_hits = {hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_661}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@221613.4]
  assign _T_668 = ~vm_enabled; // @[TLB.scala 211:18:chipyard.TestHarness.RocketConfig.fir@221614.4]
  assign hits = {_T_668,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,_T_661}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@221615.4]
  assign _GEN_33 = 2'h1 == vpn[1:0] ? sectored_entries_0_data_1 : sectored_entries_0_data_0; // @[:chipyard.TestHarness.RocketConfig.fir@221622.4]
  assign _GEN_34 = 2'h2 == vpn[1:0] ? sectored_entries_0_data_2 : _GEN_33; // @[:chipyard.TestHarness.RocketConfig.fir@221622.4]
  assign _GEN_35 = 2'h3 == vpn[1:0] ? sectored_entries_0_data_3 : _GEN_34; // @[:chipyard.TestHarness.RocketConfig.fir@221622.4]
  assign _GEN_37 = 2'h1 == vpn[1:0] ? sectored_entries_1_data_1 : sectored_entries_1_data_0; // @[:chipyard.TestHarness.RocketConfig.fir@221663.4]
  assign _GEN_38 = 2'h2 == vpn[1:0] ? sectored_entries_1_data_2 : _GEN_37; // @[:chipyard.TestHarness.RocketConfig.fir@221663.4]
  assign _GEN_39 = 2'h3 == vpn[1:0] ? sectored_entries_1_data_3 : _GEN_38; // @[:chipyard.TestHarness.RocketConfig.fir@221663.4]
  assign _GEN_41 = 2'h1 == vpn[1:0] ? sectored_entries_2_data_1 : sectored_entries_2_data_0; // @[:chipyard.TestHarness.RocketConfig.fir@221704.4]
  assign _GEN_42 = 2'h2 == vpn[1:0] ? sectored_entries_2_data_2 : _GEN_41; // @[:chipyard.TestHarness.RocketConfig.fir@221704.4]
  assign _GEN_43 = 2'h3 == vpn[1:0] ? sectored_entries_2_data_3 : _GEN_42; // @[:chipyard.TestHarness.RocketConfig.fir@221704.4]
  assign _GEN_45 = 2'h1 == vpn[1:0] ? sectored_entries_3_data_1 : sectored_entries_3_data_0; // @[:chipyard.TestHarness.RocketConfig.fir@221745.4]
  assign _GEN_46 = 2'h2 == vpn[1:0] ? sectored_entries_3_data_2 : _GEN_45; // @[:chipyard.TestHarness.RocketConfig.fir@221745.4]
  assign _GEN_47 = 2'h3 == vpn[1:0] ? sectored_entries_3_data_3 : _GEN_46; // @[:chipyard.TestHarness.RocketConfig.fir@221745.4]
  assign _GEN_49 = 2'h1 == vpn[1:0] ? sectored_entries_4_data_1 : sectored_entries_4_data_0; // @[:chipyard.TestHarness.RocketConfig.fir@221786.4]
  assign _GEN_50 = 2'h2 == vpn[1:0] ? sectored_entries_4_data_2 : _GEN_49; // @[:chipyard.TestHarness.RocketConfig.fir@221786.4]
  assign _GEN_51 = 2'h3 == vpn[1:0] ? sectored_entries_4_data_3 : _GEN_50; // @[:chipyard.TestHarness.RocketConfig.fir@221786.4]
  assign _GEN_53 = 2'h1 == vpn[1:0] ? sectored_entries_5_data_1 : sectored_entries_5_data_0; // @[:chipyard.TestHarness.RocketConfig.fir@221827.4]
  assign _GEN_54 = 2'h2 == vpn[1:0] ? sectored_entries_5_data_2 : _GEN_53; // @[:chipyard.TestHarness.RocketConfig.fir@221827.4]
  assign _GEN_55 = 2'h3 == vpn[1:0] ? sectored_entries_5_data_3 : _GEN_54; // @[:chipyard.TestHarness.RocketConfig.fir@221827.4]
  assign _GEN_57 = 2'h1 == vpn[1:0] ? sectored_entries_6_data_1 : sectored_entries_6_data_0; // @[:chipyard.TestHarness.RocketConfig.fir@221868.4]
  assign _GEN_58 = 2'h2 == vpn[1:0] ? sectored_entries_6_data_2 : _GEN_57; // @[:chipyard.TestHarness.RocketConfig.fir@221868.4]
  assign _GEN_59 = 2'h3 == vpn[1:0] ? sectored_entries_6_data_3 : _GEN_58; // @[:chipyard.TestHarness.RocketConfig.fir@221868.4]
  assign _GEN_61 = 2'h1 == vpn[1:0] ? sectored_entries_7_data_1 : sectored_entries_7_data_0; // @[:chipyard.TestHarness.RocketConfig.fir@221909.4]
  assign _GEN_62 = 2'h2 == vpn[1:0] ? sectored_entries_7_data_2 : _GEN_61; // @[:chipyard.TestHarness.RocketConfig.fir@221909.4]
  assign _GEN_63 = 2'h3 == vpn[1:0] ? sectored_entries_7_data_3 : _GEN_62; // @[:chipyard.TestHarness.RocketConfig.fir@221909.4]
  assign _T_834 = _T_439 ? vpn : 27'h0; // @[TLB.scala 108:28:chipyard.TestHarness.RocketConfig.fir@221988.4]
  assign _GEN_952 = {{7'd0}, package_Anon_9_io_y_ppn}; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@221989.4]
  assign _T_835 = _T_834 | _GEN_952; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@221989.4]
  assign _T_841 = vpn | _GEN_952; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@221995.4]
  assign _T_843 = {package_Anon_9_io_y_ppn[19:18],_T_835[17:9],_T_841[8:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@221997.4]
  assign _T_864 = _T_459 ? vpn : 27'h0; // @[TLB.scala 108:28:chipyard.TestHarness.RocketConfig.fir@222041.4]
  assign _GEN_954 = {{7'd0}, package_Anon_10_io_y_ppn}; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222042.4]
  assign _T_865 = _T_864 | _GEN_954; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222042.4]
  assign _T_871 = vpn | _GEN_954; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222048.4]
  assign _T_873 = {package_Anon_10_io_y_ppn[19:18],_T_865[17:9],_T_871[8:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@222050.4]
  assign _T_894 = _T_479 ? vpn : 27'h0; // @[TLB.scala 108:28:chipyard.TestHarness.RocketConfig.fir@222094.4]
  assign _GEN_956 = {{7'd0}, package_Anon_11_io_y_ppn}; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222095.4]
  assign _T_895 = _T_894 | _GEN_956; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222095.4]
  assign _T_901 = vpn | _GEN_956; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222101.4]
  assign _T_903 = {package_Anon_11_io_y_ppn[19:18],_T_895[17:9],_T_901[8:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@222103.4]
  assign _T_924 = _T_499 ? vpn : 27'h0; // @[TLB.scala 108:28:chipyard.TestHarness.RocketConfig.fir@222147.4]
  assign _GEN_958 = {{7'd0}, package_Anon_12_io_y_ppn}; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222148.4]
  assign _T_925 = _T_924 | _GEN_958; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222148.4]
  assign _T_931 = vpn | _GEN_958; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222154.4]
  assign _T_933 = {package_Anon_12_io_y_ppn[19:18],_T_925[17:9],_T_931[8:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@222156.4]
  assign _GEN_960 = {{7'd0}, package_Anon_13_io_y_ppn}; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222201.4]
  assign _T_955 = _T_27 | _GEN_960; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222201.4]
  assign _T_961 = _T_33 | _GEN_960; // @[TLB.scala 108:47:chipyard.TestHarness.RocketConfig.fir@222207.4]
  assign _T_963 = {package_Anon_13_io_y_ppn[19:18],_T_955[17:9],_T_961[8:0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@222209.4]
  assign _T_965 = hitsVec_0 ? package_Anon_1_io_y_ppn : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222211.4]
  assign _T_966 = hitsVec_1 ? package_Anon_2_io_y_ppn : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222212.4]
  assign _T_967 = hitsVec_2 ? package_Anon_3_io_y_ppn : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222213.4]
  assign _T_968 = hitsVec_3 ? package_Anon_4_io_y_ppn : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222214.4]
  assign _T_969 = hitsVec_4 ? package_Anon_5_io_y_ppn : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222215.4]
  assign _T_970 = hitsVec_5 ? package_Anon_6_io_y_ppn : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222216.4]
  assign _T_971 = hitsVec_6 ? package_Anon_7_io_y_ppn : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222217.4]
  assign _T_972 = hitsVec_7 ? package_Anon_8_io_y_ppn : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222218.4]
  assign _T_973 = hitsVec_8 ? _T_843 : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222219.4]
  assign _T_974 = hitsVec_9 ? _T_873 : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222220.4]
  assign _T_975 = hitsVec_10 ? _T_903 : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222221.4]
  assign _T_976 = hitsVec_11 ? _T_933 : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222222.4]
  assign _T_977 = hitsVec_12 ? _T_963 : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222223.4]
  assign _T_978 = _T_668 ? vpn[19:0] : 20'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222224.4]
  assign _T_979 = _T_965 | _T_966; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222225.4]
  assign _T_980 = _T_979 | _T_967; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222226.4]
  assign _T_981 = _T_980 | _T_968; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222227.4]
  assign _T_982 = _T_981 | _T_969; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222228.4]
  assign _T_983 = _T_982 | _T_970; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222229.4]
  assign _T_984 = _T_983 | _T_971; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222230.4]
  assign _T_985 = _T_984 | _T_972; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222231.4]
  assign _T_986 = _T_985 | _T_973; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222232.4]
  assign _T_987 = _T_986 | _T_974; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222233.4]
  assign _T_988 = _T_987 | _T_975; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222234.4]
  assign _T_989 = _T_988 | _T_976; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222235.4]
  assign _T_990 = _T_989 | _T_977; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222236.4]
  assign ppn = _T_990 | _T_978; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@222237.4]
  assign _T_992 = ~invalidate_refill; // @[TLB.scala 215:22:chipyard.TestHarness.RocketConfig.fir@222240.4]
  assign _T_993 = io_ptw_resp_valid & _T_992; // @[TLB.scala 215:19:chipyard.TestHarness.RocketConfig.fir@222241.4]
  assign _T_995 = io_ptw_resp_bits_pte_g & io_ptw_resp_bits_pte_v; // @[TLB.scala 221:25:chipyard.TestHarness.RocketConfig.fir@222248.6]
  assign _T_996 = ~io_ptw_resp_bits_pte_w; // @[PTW.scala 69:47:chipyard.TestHarness.RocketConfig.fir@222251.6]
  assign _T_997 = io_ptw_resp_bits_pte_x & _T_996; // @[PTW.scala 69:44:chipyard.TestHarness.RocketConfig.fir@222252.6]
  assign _T_998 = io_ptw_resp_bits_pte_r | _T_997; // @[PTW.scala 69:38:chipyard.TestHarness.RocketConfig.fir@222253.6]
  assign _T_999 = io_ptw_resp_bits_pte_v & _T_998; // @[PTW.scala 69:32:chipyard.TestHarness.RocketConfig.fir@222254.6]
  assign _T_1000 = _T_999 & io_ptw_resp_bits_pte_a; // @[PTW.scala 69:52:chipyard.TestHarness.RocketConfig.fir@222255.6]
  assign _T_1001 = _T_1000 & io_ptw_resp_bits_pte_r; // @[PTW.scala 73:35:chipyard.TestHarness.RocketConfig.fir@222256.6]
  assign _T_1007 = _T_1000 & io_ptw_resp_bits_pte_w; // @[PTW.scala 74:35:chipyard.TestHarness.RocketConfig.fir@222263.6]
  assign _T_1008 = _T_1007 & io_ptw_resp_bits_pte_d; // @[PTW.scala 74:40:chipyard.TestHarness.RocketConfig.fir@222264.6]
  assign _T_1014 = _T_1000 & io_ptw_resp_bits_pte_x; // @[PTW.scala 75:35:chipyard.TestHarness.RocketConfig.fir@222271.6]
  assign _T_1015 = ~io_ptw_resp_bits_homogeneous; // @[TLB.scala 234:37:chipyard.TestHarness.RocketConfig.fir@222280.6]
  assign _T_1023 = {prot_x,prot_r,_T_238,_T_238,prot_eff,cacheable,1'h0}; // @[TLB.scala 122:24:chipyard.TestHarness.RocketConfig.fir@222292.8]
  assign _T_1031 = {refill_ppn,io_ptw_resp_bits_pte_u,_T_995,io_ptw_resp_bits_ae,_T_1008,_T_1014,_T_1001,prot_w,_T_1023}; // @[TLB.scala 122:24:chipyard.TestHarness.RocketConfig.fir@222300.8]
  assign _T_1032 = io_ptw_resp_bits_level < 2'h2; // @[TLB.scala 236:40:chipyard.TestHarness.RocketConfig.fir@222304.8]
  assign _T_1033 = r_superpage_repl_addr == 2'h0; // @[TLB.scala 237:82:chipyard.TestHarness.RocketConfig.fir@222306.10]
  assign _GEN_66 = _T_1033 | superpage_entries_0_valid_0; // @[TLB.scala 237:89:chipyard.TestHarness.RocketConfig.fir@222307.10]
  assign _T_1049 = r_superpage_repl_addr == 2'h1; // @[TLB.scala 237:82:chipyard.TestHarness.RocketConfig.fir@222328.10]
  assign _GEN_70 = _T_1049 | superpage_entries_1_valid_0; // @[TLB.scala 237:89:chipyard.TestHarness.RocketConfig.fir@222329.10]
  assign _T_1065 = r_superpage_repl_addr == 2'h2; // @[TLB.scala 237:82:chipyard.TestHarness.RocketConfig.fir@222350.10]
  assign _GEN_74 = _T_1065 | superpage_entries_2_valid_0; // @[TLB.scala 237:89:chipyard.TestHarness.RocketConfig.fir@222351.10]
  assign _T_1081 = r_superpage_repl_addr == 2'h3; // @[TLB.scala 237:82:chipyard.TestHarness.RocketConfig.fir@222372.10]
  assign _GEN_78 = _T_1081 | superpage_entries_3_valid_0; // @[TLB.scala 237:89:chipyard.TestHarness.RocketConfig.fir@222373.10]
  assign _T_1097 = r_sectored_hit ? r_sectored_hit_addr : r_sectored_repl_addr; // @[TLB.scala 241:22:chipyard.TestHarness.RocketConfig.fir@222396.10]
  assign _T_1098 = _T_1097 == 3'h0; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222397.10]
  assign _T_1099 = ~r_sectored_hit; // @[TLB.scala 243:15:chipyard.TestHarness.RocketConfig.fir@222399.12]
  assign _GEN_80 = _T_1099 ? 1'h0 : sectored_entries_0_valid_0; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222400.12]
  assign _GEN_81 = _T_1099 ? 1'h0 : sectored_entries_0_valid_1; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222400.12]
  assign _GEN_82 = _T_1099 ? 1'h0 : sectored_entries_0_valid_2; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222400.12]
  assign _GEN_83 = _T_1099 ? 1'h0 : sectored_entries_0_valid_3; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222400.12]
  assign _GEN_962 = 2'h0 == r_refill_tag[1:0]; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  assign _GEN_84 = _GEN_962 | _GEN_80; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  assign _GEN_963 = 2'h1 == r_refill_tag[1:0]; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  assign _GEN_85 = _GEN_963 | _GEN_81; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  assign _GEN_964 = 2'h2 == r_refill_tag[1:0]; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  assign _GEN_86 = _GEN_964 | _GEN_82; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  assign _GEN_965 = 2'h3 == r_refill_tag[1:0]; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  assign _GEN_87 = _GEN_965 | _GEN_83; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222409.12]
  assign _GEN_92 = _T_1098 ? _GEN_84 : sectored_entries_0_valid_0; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222398.10]
  assign _GEN_93 = _T_1098 ? _GEN_85 : sectored_entries_0_valid_1; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222398.10]
  assign _GEN_94 = _T_1098 ? _GEN_86 : sectored_entries_0_valid_2; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222398.10]
  assign _GEN_95 = _T_1098 ? _GEN_87 : sectored_entries_0_valid_3; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222398.10]
  assign _T_1115 = _T_1097 == 3'h1; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222426.10]
  assign _GEN_102 = _T_1099 ? 1'h0 : sectored_entries_1_valid_0; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222429.12]
  assign _GEN_103 = _T_1099 ? 1'h0 : sectored_entries_1_valid_1; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222429.12]
  assign _GEN_104 = _T_1099 ? 1'h0 : sectored_entries_1_valid_2; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222429.12]
  assign _GEN_105 = _T_1099 ? 1'h0 : sectored_entries_1_valid_3; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222429.12]
  assign _GEN_106 = _GEN_962 | _GEN_102; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222438.12]
  assign _GEN_107 = _GEN_963 | _GEN_103; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222438.12]
  assign _GEN_108 = _GEN_964 | _GEN_104; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222438.12]
  assign _GEN_109 = _GEN_965 | _GEN_105; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222438.12]
  assign _GEN_114 = _T_1115 ? _GEN_106 : sectored_entries_1_valid_0; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222427.10]
  assign _GEN_115 = _T_1115 ? _GEN_107 : sectored_entries_1_valid_1; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222427.10]
  assign _GEN_116 = _T_1115 ? _GEN_108 : sectored_entries_1_valid_2; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222427.10]
  assign _GEN_117 = _T_1115 ? _GEN_109 : sectored_entries_1_valid_3; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222427.10]
  assign _T_1132 = _T_1097 == 3'h2; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222455.10]
  assign _GEN_124 = _T_1099 ? 1'h0 : sectored_entries_2_valid_0; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222458.12]
  assign _GEN_125 = _T_1099 ? 1'h0 : sectored_entries_2_valid_1; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222458.12]
  assign _GEN_126 = _T_1099 ? 1'h0 : sectored_entries_2_valid_2; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222458.12]
  assign _GEN_127 = _T_1099 ? 1'h0 : sectored_entries_2_valid_3; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222458.12]
  assign _GEN_128 = _GEN_962 | _GEN_124; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222467.12]
  assign _GEN_129 = _GEN_963 | _GEN_125; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222467.12]
  assign _GEN_130 = _GEN_964 | _GEN_126; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222467.12]
  assign _GEN_131 = _GEN_965 | _GEN_127; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222467.12]
  assign _GEN_136 = _T_1132 ? _GEN_128 : sectored_entries_2_valid_0; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222456.10]
  assign _GEN_137 = _T_1132 ? _GEN_129 : sectored_entries_2_valid_1; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222456.10]
  assign _GEN_138 = _T_1132 ? _GEN_130 : sectored_entries_2_valid_2; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222456.10]
  assign _GEN_139 = _T_1132 ? _GEN_131 : sectored_entries_2_valid_3; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222456.10]
  assign _T_1149 = _T_1097 == 3'h3; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222484.10]
  assign _GEN_146 = _T_1099 ? 1'h0 : sectored_entries_3_valid_0; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222487.12]
  assign _GEN_147 = _T_1099 ? 1'h0 : sectored_entries_3_valid_1; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222487.12]
  assign _GEN_148 = _T_1099 ? 1'h0 : sectored_entries_3_valid_2; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222487.12]
  assign _GEN_149 = _T_1099 ? 1'h0 : sectored_entries_3_valid_3; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222487.12]
  assign _GEN_150 = _GEN_962 | _GEN_146; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222496.12]
  assign _GEN_151 = _GEN_963 | _GEN_147; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222496.12]
  assign _GEN_152 = _GEN_964 | _GEN_148; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222496.12]
  assign _GEN_153 = _GEN_965 | _GEN_149; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222496.12]
  assign _GEN_158 = _T_1149 ? _GEN_150 : sectored_entries_3_valid_0; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222485.10]
  assign _GEN_159 = _T_1149 ? _GEN_151 : sectored_entries_3_valid_1; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222485.10]
  assign _GEN_160 = _T_1149 ? _GEN_152 : sectored_entries_3_valid_2; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222485.10]
  assign _GEN_161 = _T_1149 ? _GEN_153 : sectored_entries_3_valid_3; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222485.10]
  assign _T_1166 = _T_1097 == 3'h4; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222513.10]
  assign _GEN_168 = _T_1099 ? 1'h0 : sectored_entries_4_valid_0; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222516.12]
  assign _GEN_169 = _T_1099 ? 1'h0 : sectored_entries_4_valid_1; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222516.12]
  assign _GEN_170 = _T_1099 ? 1'h0 : sectored_entries_4_valid_2; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222516.12]
  assign _GEN_171 = _T_1099 ? 1'h0 : sectored_entries_4_valid_3; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222516.12]
  assign _GEN_172 = _GEN_962 | _GEN_168; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222525.12]
  assign _GEN_173 = _GEN_963 | _GEN_169; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222525.12]
  assign _GEN_174 = _GEN_964 | _GEN_170; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222525.12]
  assign _GEN_175 = _GEN_965 | _GEN_171; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222525.12]
  assign _GEN_180 = _T_1166 ? _GEN_172 : sectored_entries_4_valid_0; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222514.10]
  assign _GEN_181 = _T_1166 ? _GEN_173 : sectored_entries_4_valid_1; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222514.10]
  assign _GEN_182 = _T_1166 ? _GEN_174 : sectored_entries_4_valid_2; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222514.10]
  assign _GEN_183 = _T_1166 ? _GEN_175 : sectored_entries_4_valid_3; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222514.10]
  assign _T_1183 = _T_1097 == 3'h5; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222542.10]
  assign _GEN_190 = _T_1099 ? 1'h0 : sectored_entries_5_valid_0; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222545.12]
  assign _GEN_191 = _T_1099 ? 1'h0 : sectored_entries_5_valid_1; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222545.12]
  assign _GEN_192 = _T_1099 ? 1'h0 : sectored_entries_5_valid_2; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222545.12]
  assign _GEN_193 = _T_1099 ? 1'h0 : sectored_entries_5_valid_3; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222545.12]
  assign _GEN_194 = _GEN_962 | _GEN_190; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222554.12]
  assign _GEN_195 = _GEN_963 | _GEN_191; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222554.12]
  assign _GEN_196 = _GEN_964 | _GEN_192; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222554.12]
  assign _GEN_197 = _GEN_965 | _GEN_193; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222554.12]
  assign _GEN_202 = _T_1183 ? _GEN_194 : sectored_entries_5_valid_0; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222543.10]
  assign _GEN_203 = _T_1183 ? _GEN_195 : sectored_entries_5_valid_1; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222543.10]
  assign _GEN_204 = _T_1183 ? _GEN_196 : sectored_entries_5_valid_2; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222543.10]
  assign _GEN_205 = _T_1183 ? _GEN_197 : sectored_entries_5_valid_3; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222543.10]
  assign _T_1200 = _T_1097 == 3'h6; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222571.10]
  assign _GEN_212 = _T_1099 ? 1'h0 : sectored_entries_6_valid_0; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222574.12]
  assign _GEN_213 = _T_1099 ? 1'h0 : sectored_entries_6_valid_1; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222574.12]
  assign _GEN_214 = _T_1099 ? 1'h0 : sectored_entries_6_valid_2; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222574.12]
  assign _GEN_215 = _T_1099 ? 1'h0 : sectored_entries_6_valid_3; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222574.12]
  assign _GEN_216 = _GEN_962 | _GEN_212; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222583.12]
  assign _GEN_217 = _GEN_963 | _GEN_213; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222583.12]
  assign _GEN_218 = _GEN_964 | _GEN_214; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222583.12]
  assign _GEN_219 = _GEN_965 | _GEN_215; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222583.12]
  assign _GEN_224 = _T_1200 ? _GEN_216 : sectored_entries_6_valid_0; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222572.10]
  assign _GEN_225 = _T_1200 ? _GEN_217 : sectored_entries_6_valid_1; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222572.10]
  assign _GEN_226 = _T_1200 ? _GEN_218 : sectored_entries_6_valid_2; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222572.10]
  assign _GEN_227 = _T_1200 ? _GEN_219 : sectored_entries_6_valid_3; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222572.10]
  assign _T_1217 = _T_1097 == 3'h7; // @[TLB.scala 242:65:chipyard.TestHarness.RocketConfig.fir@222600.10]
  assign _GEN_234 = _T_1099 ? 1'h0 : sectored_entries_7_valid_0; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222603.12]
  assign _GEN_235 = _T_1099 ? 1'h0 : sectored_entries_7_valid_1; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222603.12]
  assign _GEN_236 = _T_1099 ? 1'h0 : sectored_entries_7_valid_2; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222603.12]
  assign _GEN_237 = _T_1099 ? 1'h0 : sectored_entries_7_valid_3; // @[TLB.scala 243:32:chipyard.TestHarness.RocketConfig.fir@222603.12]
  assign _GEN_238 = _GEN_962 | _GEN_234; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222612.12]
  assign _GEN_239 = _GEN_963 | _GEN_235; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222612.12]
  assign _GEN_240 = _GEN_964 | _GEN_236; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222612.12]
  assign _GEN_241 = _GEN_965 | _GEN_237; // @[TLB.scala 121:16:chipyard.TestHarness.RocketConfig.fir@222612.12]
  assign _GEN_246 = _T_1217 ? _GEN_238 : sectored_entries_7_valid_0; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222601.10]
  assign _GEN_247 = _T_1217 ? _GEN_239 : sectored_entries_7_valid_1; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222601.10]
  assign _GEN_248 = _T_1217 ? _GEN_240 : sectored_entries_7_valid_2; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222601.10]
  assign _GEN_249 = _T_1217 ? _GEN_241 : sectored_entries_7_valid_3; // @[TLB.scala 242:72:chipyard.TestHarness.RocketConfig.fir@222601.10]
  assign _GEN_258 = _T_1032 ? _GEN_66 : superpage_entries_0_valid_0; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_262 = _T_1032 ? _GEN_70 : superpage_entries_1_valid_0; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_266 = _T_1032 ? _GEN_74 : superpage_entries_2_valid_0; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_270 = _T_1032 ? _GEN_78 : superpage_entries_3_valid_0; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_272 = _T_1032 ? sectored_entries_0_valid_0 : _GEN_92; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_273 = _T_1032 ? sectored_entries_0_valid_1 : _GEN_93; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_274 = _T_1032 ? sectored_entries_0_valid_2 : _GEN_94; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_275 = _T_1032 ? sectored_entries_0_valid_3 : _GEN_95; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_282 = _T_1032 ? sectored_entries_1_valid_0 : _GEN_114; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_283 = _T_1032 ? sectored_entries_1_valid_1 : _GEN_115; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_284 = _T_1032 ? sectored_entries_1_valid_2 : _GEN_116; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_285 = _T_1032 ? sectored_entries_1_valid_3 : _GEN_117; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_292 = _T_1032 ? sectored_entries_2_valid_0 : _GEN_136; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_293 = _T_1032 ? sectored_entries_2_valid_1 : _GEN_137; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_294 = _T_1032 ? sectored_entries_2_valid_2 : _GEN_138; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_295 = _T_1032 ? sectored_entries_2_valid_3 : _GEN_139; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_302 = _T_1032 ? sectored_entries_3_valid_0 : _GEN_158; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_303 = _T_1032 ? sectored_entries_3_valid_1 : _GEN_159; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_304 = _T_1032 ? sectored_entries_3_valid_2 : _GEN_160; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_305 = _T_1032 ? sectored_entries_3_valid_3 : _GEN_161; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_312 = _T_1032 ? sectored_entries_4_valid_0 : _GEN_180; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_313 = _T_1032 ? sectored_entries_4_valid_1 : _GEN_181; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_314 = _T_1032 ? sectored_entries_4_valid_2 : _GEN_182; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_315 = _T_1032 ? sectored_entries_4_valid_3 : _GEN_183; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_322 = _T_1032 ? sectored_entries_5_valid_0 : _GEN_202; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_323 = _T_1032 ? sectored_entries_5_valid_1 : _GEN_203; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_324 = _T_1032 ? sectored_entries_5_valid_2 : _GEN_204; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_325 = _T_1032 ? sectored_entries_5_valid_3 : _GEN_205; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_332 = _T_1032 ? sectored_entries_6_valid_0 : _GEN_224; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_333 = _T_1032 ? sectored_entries_6_valid_1 : _GEN_225; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_334 = _T_1032 ? sectored_entries_6_valid_2 : _GEN_226; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_335 = _T_1032 ? sectored_entries_6_valid_3 : _GEN_227; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_342 = _T_1032 ? sectored_entries_7_valid_0 : _GEN_246; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_343 = _T_1032 ? sectored_entries_7_valid_1 : _GEN_247; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_344 = _T_1032 ? sectored_entries_7_valid_2 : _GEN_248; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_345 = _T_1032 ? sectored_entries_7_valid_3 : _GEN_249; // @[TLB.scala 236:54:chipyard.TestHarness.RocketConfig.fir@222305.8]
  assign _GEN_354 = _T_1015 | special_entry_valid_0; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_358 = _T_1015 ? superpage_entries_0_valid_0 : _GEN_258; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_362 = _T_1015 ? superpage_entries_1_valid_0 : _GEN_262; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_366 = _T_1015 ? superpage_entries_2_valid_0 : _GEN_266; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_370 = _T_1015 ? superpage_entries_3_valid_0 : _GEN_270; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_372 = _T_1015 ? sectored_entries_0_valid_0 : _GEN_272; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_373 = _T_1015 ? sectored_entries_0_valid_1 : _GEN_273; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_374 = _T_1015 ? sectored_entries_0_valid_2 : _GEN_274; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_375 = _T_1015 ? sectored_entries_0_valid_3 : _GEN_275; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_382 = _T_1015 ? sectored_entries_1_valid_0 : _GEN_282; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_383 = _T_1015 ? sectored_entries_1_valid_1 : _GEN_283; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_384 = _T_1015 ? sectored_entries_1_valid_2 : _GEN_284; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_385 = _T_1015 ? sectored_entries_1_valid_3 : _GEN_285; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_392 = _T_1015 ? sectored_entries_2_valid_0 : _GEN_292; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_393 = _T_1015 ? sectored_entries_2_valid_1 : _GEN_293; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_394 = _T_1015 ? sectored_entries_2_valid_2 : _GEN_294; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_395 = _T_1015 ? sectored_entries_2_valid_3 : _GEN_295; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_402 = _T_1015 ? sectored_entries_3_valid_0 : _GEN_302; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_403 = _T_1015 ? sectored_entries_3_valid_1 : _GEN_303; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_404 = _T_1015 ? sectored_entries_3_valid_2 : _GEN_304; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_405 = _T_1015 ? sectored_entries_3_valid_3 : _GEN_305; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_412 = _T_1015 ? sectored_entries_4_valid_0 : _GEN_312; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_413 = _T_1015 ? sectored_entries_4_valid_1 : _GEN_313; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_414 = _T_1015 ? sectored_entries_4_valid_2 : _GEN_314; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_415 = _T_1015 ? sectored_entries_4_valid_3 : _GEN_315; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_422 = _T_1015 ? sectored_entries_5_valid_0 : _GEN_322; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_423 = _T_1015 ? sectored_entries_5_valid_1 : _GEN_323; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_424 = _T_1015 ? sectored_entries_5_valid_2 : _GEN_324; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_425 = _T_1015 ? sectored_entries_5_valid_3 : _GEN_325; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_432 = _T_1015 ? sectored_entries_6_valid_0 : _GEN_332; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_433 = _T_1015 ? sectored_entries_6_valid_1 : _GEN_333; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_434 = _T_1015 ? sectored_entries_6_valid_2 : _GEN_334; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_435 = _T_1015 ? sectored_entries_6_valid_3 : _GEN_335; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_442 = _T_1015 ? sectored_entries_7_valid_0 : _GEN_342; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_443 = _T_1015 ? sectored_entries_7_valid_1 : _GEN_343; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_444 = _T_1015 ? sectored_entries_7_valid_2 : _GEN_344; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_445 = _T_1015 ? sectored_entries_7_valid_3 : _GEN_345; // @[TLB.scala 234:68:chipyard.TestHarness.RocketConfig.fir@222282.6]
  assign _GEN_454 = _T_993 ? _GEN_354 : special_entry_valid_0; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_458 = _T_993 ? _GEN_358 : superpage_entries_0_valid_0; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_462 = _T_993 ? _GEN_362 : superpage_entries_1_valid_0; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_466 = _T_993 ? _GEN_366 : superpage_entries_2_valid_0; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_470 = _T_993 ? _GEN_370 : superpage_entries_3_valid_0; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_472 = _T_993 ? _GEN_372 : sectored_entries_0_valid_0; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_473 = _T_993 ? _GEN_373 : sectored_entries_0_valid_1; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_474 = _T_993 ? _GEN_374 : sectored_entries_0_valid_2; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_475 = _T_993 ? _GEN_375 : sectored_entries_0_valid_3; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_482 = _T_993 ? _GEN_382 : sectored_entries_1_valid_0; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_483 = _T_993 ? _GEN_383 : sectored_entries_1_valid_1; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_484 = _T_993 ? _GEN_384 : sectored_entries_1_valid_2; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_485 = _T_993 ? _GEN_385 : sectored_entries_1_valid_3; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_492 = _T_993 ? _GEN_392 : sectored_entries_2_valid_0; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_493 = _T_993 ? _GEN_393 : sectored_entries_2_valid_1; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_494 = _T_993 ? _GEN_394 : sectored_entries_2_valid_2; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_495 = _T_993 ? _GEN_395 : sectored_entries_2_valid_3; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_502 = _T_993 ? _GEN_402 : sectored_entries_3_valid_0; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_503 = _T_993 ? _GEN_403 : sectored_entries_3_valid_1; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_504 = _T_993 ? _GEN_404 : sectored_entries_3_valid_2; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_505 = _T_993 ? _GEN_405 : sectored_entries_3_valid_3; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_512 = _T_993 ? _GEN_412 : sectored_entries_4_valid_0; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_513 = _T_993 ? _GEN_413 : sectored_entries_4_valid_1; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_514 = _T_993 ? _GEN_414 : sectored_entries_4_valid_2; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_515 = _T_993 ? _GEN_415 : sectored_entries_4_valid_3; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_522 = _T_993 ? _GEN_422 : sectored_entries_5_valid_0; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_523 = _T_993 ? _GEN_423 : sectored_entries_5_valid_1; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_524 = _T_993 ? _GEN_424 : sectored_entries_5_valid_2; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_525 = _T_993 ? _GEN_425 : sectored_entries_5_valid_3; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_532 = _T_993 ? _GEN_432 : sectored_entries_6_valid_0; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_533 = _T_993 ? _GEN_433 : sectored_entries_6_valid_1; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_534 = _T_993 ? _GEN_434 : sectored_entries_6_valid_2; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_535 = _T_993 ? _GEN_435 : sectored_entries_6_valid_3; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_542 = _T_993 ? _GEN_442 : sectored_entries_7_valid_0; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_543 = _T_993 ? _GEN_443 : sectored_entries_7_valid_1; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_544 = _T_993 ? _GEN_444 : sectored_entries_7_valid_2; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _GEN_545 = _T_993 ? _GEN_445 : sectored_entries_7_valid_3; // @[TLB.scala 215:42:chipyard.TestHarness.RocketConfig.fir@222242.4]
  assign _T_1679 = {package_Anon_19_io_y_ae,package_Anon_18_io_y_ae,package_Anon_17_io_y_ae,package_Anon_16_io_y_ae,package_Anon_15_io_y_ae,package_Anon_14_io_y_ae}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223651.4]
  assign ptw_ae_array = {1'h0,package_Anon_26_io_y_ae,package_Anon_25_io_y_ae,package_Anon_24_io_y_ae,package_Anon_23_io_y_ae,package_Anon_22_io_y_ae,package_Anon_21_io_y_ae,package_Anon_20_io_y_ae,_T_1679}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223659.4]
  assign _T_1693 = {package_Anon_19_io_y_u,package_Anon_18_io_y_u,package_Anon_17_io_y_u,package_Anon_16_io_y_u,package_Anon_15_io_y_u,package_Anon_14_io_y_u}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223666.4]
  assign _T_1700 = {package_Anon_26_io_y_u,package_Anon_25_io_y_u,package_Anon_24_io_y_u,package_Anon_23_io_y_u,package_Anon_22_io_y_u,package_Anon_21_io_y_u,package_Anon_20_io_y_u,_T_1693}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223673.4]
  assign _T_1714 = ~_T_1700; // @[TLB.scala 253:98:chipyard.TestHarness.RocketConfig.fir@223687.4]
  assign priv_x_ok = priv_s ? _T_1714 : _T_1700; // @[TLB.scala 254:22:chipyard.TestHarness.RocketConfig.fir@223715.4]
  assign _T_1757 = {package_Anon_19_io_y_sx,package_Anon_18_io_y_sx,package_Anon_17_io_y_sx,package_Anon_16_io_y_sx,package_Anon_15_io_y_sx,package_Anon_14_io_y_sx}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223732.4]
  assign _T_1764 = {package_Anon_26_io_y_sx,package_Anon_25_io_y_sx,package_Anon_24_io_y_sx,package_Anon_23_io_y_sx,package_Anon_22_io_y_sx,package_Anon_21_io_y_sx,package_Anon_20_io_y_sx,_T_1757}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223739.4]
  assign _T_1793 = priv_x_ok & _T_1764; // @[TLB.scala 257:39:chipyard.TestHarness.RocketConfig.fir@223770.4]
  assign x_array = {1'h1,_T_1793}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223771.4]
  assign _T_1808 = ~ptw_ae_array; // @[TLB.scala 258:89:chipyard.TestHarness.RocketConfig.fir@223786.4]
  assign _T_1825 = prot_x ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@223805.4]
  assign _T_1830 = {package_Anon_32_io_y_px,package_Anon_31_io_y_px,package_Anon_30_io_y_px,package_Anon_29_io_y_px,package_Anon_28_io_y_px,package_Anon_27_io_y_px}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223810.4]
  assign _T_1837 = {_T_1825,package_Anon_38_io_y_px,package_Anon_37_io_y_px,package_Anon_36_io_y_px,package_Anon_35_io_y_px,package_Anon_34_io_y_px,package_Anon_33_io_y_px,_T_1830}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223817.4]
  assign px_array = _T_1837 & _T_1808; // @[TLB.scala 260:87:chipyard.TestHarness.RocketConfig.fir@223819.4]
  assign _T_1853 = cacheable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@223835.4]
  assign _T_1858 = {package_Anon_32_io_y_c,package_Anon_31_io_y_c,package_Anon_30_io_y_c,package_Anon_29_io_y_c,package_Anon_28_io_y_c,package_Anon_27_io_y_c}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223840.4]
  assign c_array = {_T_1853,package_Anon_38_io_y_c,package_Anon_37_io_y_c,package_Anon_36_io_y_c,package_Anon_35_io_y_c,package_Anon_34_io_y_c,package_Anon_33_io_y_c,_T_1858}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@223847.4]
  assign _T_1910 = io_req_bits_vaddr & 40'hc000000000; // @[TLB.scala 275:43:chipyard.TestHarness.RocketConfig.fir@223899.4]
  assign _T_1912 = _T_1910 == 40'h0; // @[TLB.scala 276:61:chipyard.TestHarness.RocketConfig.fir@223901.4]
  assign _T_1913 = _T_1910 == 40'hc000000000; // @[TLB.scala 276:82:chipyard.TestHarness.RocketConfig.fir@223902.4]
  assign _T_1914 = _T_1912 | _T_1913; // @[TLB.scala 276:67:chipyard.TestHarness.RocketConfig.fir@223903.4]
  assign _T_1915 = ~_T_1914; // @[TLB.scala 276:47:chipyard.TestHarness.RocketConfig.fir@223904.4]
  assign bad_va = vm_enabled & _T_1915; // @[TLB.scala 270:117:chipyard.TestHarness.RocketConfig.fir@223906.4]
  assign _T_2011 = x_array | ptw_ae_array; // @[TLB.scala 305:33:chipyard.TestHarness.RocketConfig.fir@224016.4]
  assign pf_inst_array = ~_T_2011; // @[TLB.scala 305:23:chipyard.TestHarness.RocketConfig.fir@224017.4]
  assign tlb_hit = |real_hits; // @[TLB.scala 307:27:chipyard.TestHarness.RocketConfig.fir@224018.4]
  assign _T_2012 = ~bad_va; // @[TLB.scala 308:32:chipyard.TestHarness.RocketConfig.fir@224019.4]
  assign _T_2013 = vm_enabled & _T_2012; // @[TLB.scala 308:29:chipyard.TestHarness.RocketConfig.fir@224020.4]
  assign _T_2014 = ~tlb_hit; // @[TLB.scala 308:43:chipyard.TestHarness.RocketConfig.fir@224021.4]
  assign tlb_miss = _T_2013 & _T_2014; // @[TLB.scala 308:40:chipyard.TestHarness.RocketConfig.fir@224022.4]
  assign _T_2017 = io_req_valid & vm_enabled; // @[TLB.scala 312:22:chipyard.TestHarness.RocketConfig.fir@224025.4]
  assign _T_2018 = sector_hits_0 | sector_hits_1; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224027.6]
  assign _T_2019 = _T_2018 | sector_hits_2; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224028.6]
  assign _T_2020 = _T_2019 | sector_hits_3; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224029.6]
  assign _T_2021 = _T_2020 | sector_hits_4; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224030.6]
  assign _T_2022 = _T_2021 | sector_hits_5; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224031.6]
  assign _T_2023 = _T_2022 | sector_hits_6; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224032.6]
  assign _T_2024 = _T_2023 | sector_hits_7; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224033.6]
  assign _T_2031 = {sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,sector_hits_0}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224041.8]
  assign _T_2034 = |_T_2031[7:4]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@224044.8]
  assign _T_2035 = _T_2031[7:4] | _T_2031[3:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@224045.8]
  assign _T_2038 = |_T_2035[3:2]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@224048.8]
  assign _T_2039 = _T_2035[3:2] | _T_2035[1:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@224049.8]
  assign _T_2042 = {_T_2034,_T_2038,_T_2039[1]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224052.8]
  assign _T_2043 = {_T_2015, 1'h0}; // @[Replacement.scala 50:28:chipyard.TestHarness.RocketConfig.fir@224053.8]
  assign _T_2045 = ~_T_2042[2]; // @[Replacement.scala 54:43:chipyard.TestHarness.RocketConfig.fir@224055.8]
  assign _T_2047 = _T_2043 | 8'h2; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224057.8]
  assign _T_2048 = ~_T_2043; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224058.8]
  assign _T_2049 = _T_2048 | 8'h2; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224059.8]
  assign _T_2050 = ~_T_2049; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224060.8]
  assign _T_2051 = _T_2045 ? _T_2047 : _T_2050; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224061.8]
  assign _T_2052 = {1'h1,_T_2042[2]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224062.8]
  assign _T_2054 = ~_T_2042[1]; // @[Replacement.scala 54:43:chipyard.TestHarness.RocketConfig.fir@224064.8]
  assign _T_2055 = 4'h1 << _T_2052; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224065.8]
  assign _GEN_995 = {{4'd0}, _T_2055}; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224066.8]
  assign _T_2056 = _T_2051 | _GEN_995; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224066.8]
  assign _T_2057 = ~_T_2051; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224067.8]
  assign _T_2058 = _T_2057 | _GEN_995; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224068.8]
  assign _T_2059 = ~_T_2058; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224069.8]
  assign _T_2060 = _T_2054 ? _T_2056 : _T_2059; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224070.8]
  assign _T_2061 = {1'h1,_T_2042[2],_T_2042[1]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224071.8]
  assign _T_2063 = ~_T_2042[0]; // @[Replacement.scala 54:43:chipyard.TestHarness.RocketConfig.fir@224073.8]
  assign _T_2064 = 8'h1 << _T_2061; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224074.8]
  assign _T_2065 = _T_2060 | _T_2064; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224075.8]
  assign _T_2066 = ~_T_2060; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224076.8]
  assign _T_2067 = _T_2066 | _T_2064; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224077.8]
  assign _T_2068 = ~_T_2067; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224078.8]
  assign _T_2069 = _T_2063 ? _T_2065 : _T_2068; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224079.8]
  assign _T_2072 = superpage_hits_0 | superpage_hits_1; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224084.6]
  assign _T_2073 = _T_2072 | superpage_hits_2; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224085.6]
  assign _T_2074 = _T_2073 | superpage_hits_3; // @[package.scala 64:59:chipyard.TestHarness.RocketConfig.fir@224086.6]
  assign _T_2077 = {superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224090.8]
  assign _T_2080 = |_T_2077[3:2]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@224093.8]
  assign _T_2081 = _T_2077[3:2] | _T_2077[1:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@224094.8]
  assign _T_2083 = {_T_2080,_T_2081[1]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224096.8]
  assign _T_2084 = {_T_2016, 1'h0}; // @[Replacement.scala 50:28:chipyard.TestHarness.RocketConfig.fir@224097.8]
  assign _T_2086 = ~_T_2083[1]; // @[Replacement.scala 54:43:chipyard.TestHarness.RocketConfig.fir@224099.8]
  assign _T_2088 = _T_2084 | 4'h2; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224101.8]
  assign _T_2089 = ~_T_2084; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224102.8]
  assign _T_2090 = _T_2089 | 4'h2; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224103.8]
  assign _T_2091 = ~_T_2090; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224104.8]
  assign _T_2092 = _T_2086 ? _T_2088 : _T_2091; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224105.8]
  assign _T_2093 = {1'h1,_T_2083[1]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224106.8]
  assign _T_2095 = ~_T_2083[0]; // @[Replacement.scala 54:43:chipyard.TestHarness.RocketConfig.fir@224108.8]
  assign _T_2096 = 4'h1 << _T_2093; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224109.8]
  assign _T_2097 = _T_2092 | _T_2096; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224110.8]
  assign _T_2098 = ~_T_2092; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224111.8]
  assign _T_2099 = _T_2098 | _T_2096; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224112.8]
  assign _T_2100 = ~_T_2099; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224113.8]
  assign _T_2101 = _T_2095 ? _T_2097 : _T_2100; // @[Replacement.scala 54:37:chipyard.TestHarness.RocketConfig.fir@224114.8]
  assign _T_2113 = real_hits[1] | real_hits[2]; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224129.4]
  assign _T_2115 = real_hits[1] & real_hits[2]; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224131.4]
  assign _T_2117 = real_hits[0] | _T_2113; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224133.4]
  assign _T_2119 = real_hits[0] & _T_2113; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224135.4]
  assign _T_2120 = _T_2115 | _T_2119; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224136.4]
  assign _T_2129 = real_hits[4] | real_hits[5]; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224145.4]
  assign _T_2131 = real_hits[4] & real_hits[5]; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224147.4]
  assign _T_2133 = real_hits[3] | _T_2129; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224149.4]
  assign _T_2135 = real_hits[3] & _T_2129; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224151.4]
  assign _T_2136 = _T_2131 | _T_2135; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224152.4]
  assign _T_2137 = _T_2117 | _T_2133; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224153.4]
  assign _T_2138 = _T_2120 | _T_2136; // @[Misc.scala 182:37:chipyard.TestHarness.RocketConfig.fir@224154.4]
  assign _T_2139 = _T_2117 & _T_2133; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224155.4]
  assign _T_2140 = _T_2138 | _T_2139; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224156.4]
  assign _T_2150 = real_hits[7] | real_hits[8]; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224166.4]
  assign _T_2152 = real_hits[7] & real_hits[8]; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224168.4]
  assign _T_2154 = real_hits[6] | _T_2150; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224170.4]
  assign _T_2156 = real_hits[6] & _T_2150; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224172.4]
  assign _T_2157 = _T_2152 | _T_2156; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224173.4]
  assign _T_2164 = real_hits[9] | real_hits[10]; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224180.4]
  assign _T_2166 = real_hits[9] & real_hits[10]; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224182.4]
  assign _T_2173 = real_hits[11] | real_hits[12]; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224189.4]
  assign _T_2175 = real_hits[11] & real_hits[12]; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224191.4]
  assign _T_2177 = _T_2164 | _T_2173; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224193.4]
  assign _T_2178 = _T_2166 | _T_2175; // @[Misc.scala 182:37:chipyard.TestHarness.RocketConfig.fir@224194.4]
  assign _T_2179 = _T_2164 & _T_2173; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224195.4]
  assign _T_2180 = _T_2178 | _T_2179; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224196.4]
  assign _T_2181 = _T_2154 | _T_2177; // @[Misc.scala 182:16:chipyard.TestHarness.RocketConfig.fir@224197.4]
  assign _T_2182 = _T_2157 | _T_2180; // @[Misc.scala 182:37:chipyard.TestHarness.RocketConfig.fir@224198.4]
  assign _T_2183 = _T_2154 & _T_2177; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224199.4]
  assign _T_2184 = _T_2182 | _T_2183; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224200.4]
  assign _T_2186 = _T_2140 | _T_2184; // @[Misc.scala 182:37:chipyard.TestHarness.RocketConfig.fir@224202.4]
  assign _T_2187 = _T_2137 & _T_2181; // @[Misc.scala 182:61:chipyard.TestHarness.RocketConfig.fir@224203.4]
  assign multipleHits = _T_2186 | _T_2187; // @[Misc.scala 182:49:chipyard.TestHarness.RocketConfig.fir@224204.4]
  assign _T_2197 = pf_inst_array & hits; // @[TLB.scala 327:47:chipyard.TestHarness.RocketConfig.fir@224217.4]
  assign _T_2198 = |_T_2197; // @[TLB.scala 327:55:chipyard.TestHarness.RocketConfig.fir@224218.4]
  assign _T_2204 = ~px_array; // @[TLB.scala 330:23:chipyard.TestHarness.RocketConfig.fir@224227.4]
  assign _T_2205 = _T_2204 & hits; // @[TLB.scala 330:33:chipyard.TestHarness.RocketConfig.fir@224228.4]
  assign _T_2211 = c_array & hits; // @[TLB.scala 334:33:chipyard.TestHarness.RocketConfig.fir@224238.4]
  assign _T_2218 = io_ptw_resp_valid | tlb_miss; // @[TLB.scala 337:29:chipyard.TestHarness.RocketConfig.fir@224248.4]
  assign _T_2224 = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37:chipyard.TestHarness.RocketConfig.fir@224259.4]
  assign _T_2225 = _T_2224 & tlb_miss; // @[TLB.scala 346:25:chipyard.TestHarness.RocketConfig.fir@224260.4]
  assign _T_2230 = {{1'd0}, _T_2084[3:1]}; // @[Replacement.scala 65:48:chipyard.TestHarness.RocketConfig.fir@224268.6]
  assign _T_2233 = {1'h1,_T_2230[0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224271.6]
  assign _T_2237 = _T_2084 >> _T_2233; // @[Replacement.scala 65:48:chipyard.TestHarness.RocketConfig.fir@224275.6]
  assign _T_2240 = {1'h1,_T_2230[0],_T_2237[0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224278.6]
  assign _T_2244 = {superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,superpage_entries_0_valid_0}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224282.6]
  assign _T_2245 = &_T_2244; // @[TLB.scala 394:16:chipyard.TestHarness.RocketConfig.fir@224283.6]
  assign _T_2246 = ~_T_2244; // @[TLB.scala 394:43:chipyard.TestHarness.RocketConfig.fir@224284.6]
  assign _T_2259 = {{1'd0}, _T_2043[7:1]}; // @[Replacement.scala 65:48:chipyard.TestHarness.RocketConfig.fir@224298.6]
  assign _T_2262 = {1'h1,_T_2259[0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224301.6]
  assign _T_2266 = _T_2043 >> _T_2262; // @[Replacement.scala 65:48:chipyard.TestHarness.RocketConfig.fir@224305.6]
  assign _T_2269 = {1'h1,_T_2259[0],_T_2266[0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224308.6]
  assign _T_2273 = _T_2043 >> _T_2269; // @[Replacement.scala 65:48:chipyard.TestHarness.RocketConfig.fir@224312.6]
  assign _T_2276 = {1'h1,_T_2259[0],_T_2266[0],_T_2273[0]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224315.6]
  assign _T_2308 = {_T_428,_T_422,_T_416,_T_410,_T_404,_T_398,_T_392,_T_386}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@224347.6]
  assign _T_2309 = &_T_2308; // @[TLB.scala 394:16:chipyard.TestHarness.RocketConfig.fir@224348.6]
  assign _T_2310 = ~_T_2308; // @[TLB.scala 394:43:chipyard.TestHarness.RocketConfig.fir@224349.6]
  assign _T_2354 = state == 2'h2; // @[TLB.scala 360:17:chipyard.TestHarness.RocketConfig.fir@224408.4]
  assign _T_2355 = _T_2354 & io_sfence_valid; // @[TLB.scala 360:28:chipyard.TestHarness.RocketConfig.fir@224409.4]
  assign _T_2356 = ~io_sfence_bits_rs1; // @[TLB.scala 368:14:chipyard.TestHarness.RocketConfig.fir@224417.6]
  assign _T_2358 = io_sfence_bits_addr[38:12] == vpn; // @[TLB.scala 368:72:chipyard.TestHarness.RocketConfig.fir@224419.6]
  assign _T_2359 = _T_2356 | _T_2358; // @[TLB.scala 368:34:chipyard.TestHarness.RocketConfig.fir@224420.6]
  assign _T_2361 = _T_2359 | reset; // @[TLB.scala 368:13:chipyard.TestHarness.RocketConfig.fir@224422.6]
  assign _T_2362 = ~_T_2361; // @[TLB.scala 368:13:chipyard.TestHarness.RocketConfig.fir@224423.6]
  assign _T_2369 = _T_387[26:18] == 9'h0; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@224438.8]
  assign _T_2506 = ~sectored_entries_0_data_0[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@224736.10]
  assign _GEN_648 = _T_2506 ? 1'h0 : _GEN_472; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@224737.10]
  assign _T_2507 = ~sectored_entries_0_data_1[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@224740.10]
  assign _GEN_649 = _T_2507 ? 1'h0 : _GEN_473; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@224741.10]
  assign _T_2508 = ~sectored_entries_0_data_2[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@224744.10]
  assign _GEN_650 = _T_2508 ? 1'h0 : _GEN_474; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@224745.10]
  assign _T_2509 = ~sectored_entries_0_data_3[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@224748.10]
  assign _GEN_651 = _T_2509 ? 1'h0 : _GEN_475; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@224749.10]
  assign _GEN_652 = io_sfence_bits_rs2 & _GEN_648; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224595.8]
  assign _GEN_653 = io_sfence_bits_rs2 & _GEN_649; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224595.8]
  assign _GEN_654 = io_sfence_bits_rs2 & _GEN_650; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224595.8]
  assign _GEN_655 = io_sfence_bits_rs2 & _GEN_651; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224595.8]
  assign _T_2516 = _T_393[26:18] == 9'h0; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@224769.8]
  assign _T_2653 = ~sectored_entries_1_data_0[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225067.10]
  assign _GEN_676 = _T_2653 ? 1'h0 : _GEN_482; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225068.10]
  assign _T_2654 = ~sectored_entries_1_data_1[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225071.10]
  assign _GEN_677 = _T_2654 ? 1'h0 : _GEN_483; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225072.10]
  assign _T_2655 = ~sectored_entries_1_data_2[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225075.10]
  assign _GEN_678 = _T_2655 ? 1'h0 : _GEN_484; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225076.10]
  assign _T_2656 = ~sectored_entries_1_data_3[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225079.10]
  assign _GEN_679 = _T_2656 ? 1'h0 : _GEN_485; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225080.10]
  assign _GEN_680 = io_sfence_bits_rs2 & _GEN_676; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224926.8]
  assign _GEN_681 = io_sfence_bits_rs2 & _GEN_677; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224926.8]
  assign _GEN_682 = io_sfence_bits_rs2 & _GEN_678; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224926.8]
  assign _GEN_683 = io_sfence_bits_rs2 & _GEN_679; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@224926.8]
  assign _T_2663 = _T_399[26:18] == 9'h0; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@225100.8]
  assign _T_2800 = ~sectored_entries_2_data_0[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225398.10]
  assign _GEN_704 = _T_2800 ? 1'h0 : _GEN_492; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225399.10]
  assign _T_2801 = ~sectored_entries_2_data_1[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225402.10]
  assign _GEN_705 = _T_2801 ? 1'h0 : _GEN_493; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225403.10]
  assign _T_2802 = ~sectored_entries_2_data_2[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225406.10]
  assign _GEN_706 = _T_2802 ? 1'h0 : _GEN_494; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225407.10]
  assign _T_2803 = ~sectored_entries_2_data_3[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225410.10]
  assign _GEN_707 = _T_2803 ? 1'h0 : _GEN_495; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225411.10]
  assign _GEN_708 = io_sfence_bits_rs2 & _GEN_704; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225257.8]
  assign _GEN_709 = io_sfence_bits_rs2 & _GEN_705; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225257.8]
  assign _GEN_710 = io_sfence_bits_rs2 & _GEN_706; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225257.8]
  assign _GEN_711 = io_sfence_bits_rs2 & _GEN_707; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225257.8]
  assign _T_2810 = _T_405[26:18] == 9'h0; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@225431.8]
  assign _T_2947 = ~sectored_entries_3_data_0[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225729.10]
  assign _GEN_732 = _T_2947 ? 1'h0 : _GEN_502; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225730.10]
  assign _T_2948 = ~sectored_entries_3_data_1[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225733.10]
  assign _GEN_733 = _T_2948 ? 1'h0 : _GEN_503; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225734.10]
  assign _T_2949 = ~sectored_entries_3_data_2[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225737.10]
  assign _GEN_734 = _T_2949 ? 1'h0 : _GEN_504; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225738.10]
  assign _T_2950 = ~sectored_entries_3_data_3[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@225741.10]
  assign _GEN_735 = _T_2950 ? 1'h0 : _GEN_505; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@225742.10]
  assign _GEN_736 = io_sfence_bits_rs2 & _GEN_732; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225588.8]
  assign _GEN_737 = io_sfence_bits_rs2 & _GEN_733; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225588.8]
  assign _GEN_738 = io_sfence_bits_rs2 & _GEN_734; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225588.8]
  assign _GEN_739 = io_sfence_bits_rs2 & _GEN_735; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225588.8]
  assign _T_2957 = _T_411[26:18] == 9'h0; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@225762.8]
  assign _T_3094 = ~sectored_entries_4_data_0[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226060.10]
  assign _GEN_760 = _T_3094 ? 1'h0 : _GEN_512; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226061.10]
  assign _T_3095 = ~sectored_entries_4_data_1[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226064.10]
  assign _GEN_761 = _T_3095 ? 1'h0 : _GEN_513; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226065.10]
  assign _T_3096 = ~sectored_entries_4_data_2[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226068.10]
  assign _GEN_762 = _T_3096 ? 1'h0 : _GEN_514; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226069.10]
  assign _T_3097 = ~sectored_entries_4_data_3[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226072.10]
  assign _GEN_763 = _T_3097 ? 1'h0 : _GEN_515; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226073.10]
  assign _GEN_764 = io_sfence_bits_rs2 & _GEN_760; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225919.8]
  assign _GEN_765 = io_sfence_bits_rs2 & _GEN_761; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225919.8]
  assign _GEN_766 = io_sfence_bits_rs2 & _GEN_762; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225919.8]
  assign _GEN_767 = io_sfence_bits_rs2 & _GEN_763; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@225919.8]
  assign _T_3104 = _T_417[26:18] == 9'h0; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@226093.8]
  assign _T_3241 = ~sectored_entries_5_data_0[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226391.10]
  assign _GEN_788 = _T_3241 ? 1'h0 : _GEN_522; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226392.10]
  assign _T_3242 = ~sectored_entries_5_data_1[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226395.10]
  assign _GEN_789 = _T_3242 ? 1'h0 : _GEN_523; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226396.10]
  assign _T_3243 = ~sectored_entries_5_data_2[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226399.10]
  assign _GEN_790 = _T_3243 ? 1'h0 : _GEN_524; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226400.10]
  assign _T_3244 = ~sectored_entries_5_data_3[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226403.10]
  assign _GEN_791 = _T_3244 ? 1'h0 : _GEN_525; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226404.10]
  assign _GEN_792 = io_sfence_bits_rs2 & _GEN_788; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226250.8]
  assign _GEN_793 = io_sfence_bits_rs2 & _GEN_789; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226250.8]
  assign _GEN_794 = io_sfence_bits_rs2 & _GEN_790; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226250.8]
  assign _GEN_795 = io_sfence_bits_rs2 & _GEN_791; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226250.8]
  assign _T_3251 = _T_423[26:18] == 9'h0; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@226424.8]
  assign _T_3388 = ~sectored_entries_6_data_0[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226722.10]
  assign _GEN_816 = _T_3388 ? 1'h0 : _GEN_532; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226723.10]
  assign _T_3389 = ~sectored_entries_6_data_1[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226726.10]
  assign _GEN_817 = _T_3389 ? 1'h0 : _GEN_533; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226727.10]
  assign _T_3390 = ~sectored_entries_6_data_2[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226730.10]
  assign _GEN_818 = _T_3390 ? 1'h0 : _GEN_534; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226731.10]
  assign _T_3391 = ~sectored_entries_6_data_3[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@226734.10]
  assign _GEN_819 = _T_3391 ? 1'h0 : _GEN_535; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@226735.10]
  assign _GEN_820 = io_sfence_bits_rs2 & _GEN_816; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226581.8]
  assign _GEN_821 = io_sfence_bits_rs2 & _GEN_817; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226581.8]
  assign _GEN_822 = io_sfence_bits_rs2 & _GEN_818; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226581.8]
  assign _GEN_823 = io_sfence_bits_rs2 & _GEN_819; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226581.8]
  assign _T_3398 = _T_429[26:18] == 9'h0; // @[TLB.scala 134:61:chipyard.TestHarness.RocketConfig.fir@226755.8]
  assign _T_3535 = ~sectored_entries_7_data_0[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227053.10]
  assign _GEN_844 = _T_3535 ? 1'h0 : _GEN_542; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227054.10]
  assign _T_3536 = ~sectored_entries_7_data_1[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227057.10]
  assign _GEN_845 = _T_3536 ? 1'h0 : _GEN_543; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227058.10]
  assign _T_3537 = ~sectored_entries_7_data_2[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227061.10]
  assign _GEN_846 = _T_3537 ? 1'h0 : _GEN_544; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227062.10]
  assign _T_3538 = ~sectored_entries_7_data_3[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227065.10]
  assign _GEN_847 = _T_3538 ? 1'h0 : _GEN_545; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227066.10]
  assign _GEN_848 = io_sfence_bits_rs2 & _GEN_844; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226912.8]
  assign _GEN_849 = io_sfence_bits_rs2 & _GEN_845; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226912.8]
  assign _GEN_850 = io_sfence_bits_rs2 & _GEN_846; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226912.8]
  assign _GEN_851 = io_sfence_bits_rs2 & _GEN_847; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@226912.8]
  assign _T_3577 = ~superpage_entries_0_data_0[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227139.10]
  assign _GEN_857 = _T_3577 ? 1'h0 : _GEN_458; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227140.10]
  assign _GEN_858 = io_sfence_bits_rs2 & _GEN_857; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@227103.8]
  assign _T_3616 = ~superpage_entries_1_data_0[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227210.10]
  assign _GEN_861 = _T_3616 ? 1'h0 : _GEN_462; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227211.10]
  assign _GEN_862 = io_sfence_bits_rs2 & _GEN_861; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@227174.8]
  assign _T_3655 = ~superpage_entries_2_data_0[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227281.10]
  assign _GEN_865 = _T_3655 ? 1'h0 : _GEN_466; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227282.10]
  assign _GEN_866 = io_sfence_bits_rs2 & _GEN_865; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@227245.8]
  assign _T_3694 = ~superpage_entries_3_data_0[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227352.10]
  assign _GEN_869 = _T_3694 ? 1'h0 : _GEN_470; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227353.10]
  assign _GEN_870 = io_sfence_bits_rs2 & _GEN_869; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@227316.8]
  assign _T_3733 = ~special_entry_data_0[12]; // @[TLB.scala 142:13:chipyard.TestHarness.RocketConfig.fir@227423.10]
  assign _GEN_873 = _T_3733 ? 1'h0 : _GEN_454; // @[TLB.scala 142:19:chipyard.TestHarness.RocketConfig.fir@227424.10]
  assign _GEN_874 = io_sfence_bits_rs2 & _GEN_873; // @[TLB.scala 371:40:chipyard.TestHarness.RocketConfig.fir@227387.8]
  assign _T_3735 = multipleHits | reset; // @[TLB.scala 375:24:chipyard.TestHarness.RocketConfig.fir@227433.4]
  assign io_req_ready = state == 2'h0; // @[TLB.scala 324:16:chipyard.TestHarness.RocketConfig.fir@224206.4]
  assign io_resp_miss = _T_2218 | multipleHits; // @[TLB.scala 337:16:chipyard.TestHarness.RocketConfig.fir@224250.4]
  assign io_resp_paddr = {ppn,io_req_bits_vaddr[11:0]}; // @[TLB.scala 338:17:chipyard.TestHarness.RocketConfig.fir@224253.4]
  assign io_resp_pf_inst = bad_va | _T_2198; // @[TLB.scala 327:19:chipyard.TestHarness.RocketConfig.fir@224220.4]
  assign io_resp_ae_inst = |_T_2205; // @[TLB.scala 330:19:chipyard.TestHarness.RocketConfig.fir@224230.4]
  assign io_resp_cacheable = |_T_2211; // @[TLB.scala 334:21:chipyard.TestHarness.RocketConfig.fir@224240.4]
  assign io_ptw_req_valid = state == 2'h1; // @[TLB.scala 340:20:chipyard.TestHarness.RocketConfig.fir@224255.4]
  assign io_ptw_req_bits_valid = ~io_kill; // @[TLB.scala 341:25:chipyard.TestHarness.RocketConfig.fir@224257.4]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[TLB.scala 342:29:chipyard.TestHarness.RocketConfig.fir@224258.4]
  assign package_Anon_io_x_ppn = special_entry_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@220900.4]
  assign package_Anon_io_x_u = special_entry_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@220900.4]
  assign package_Anon_io_x_ae = special_entry_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@220900.4]
  assign package_Anon_io_x_sw = special_entry_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@220900.4]
  assign package_Anon_io_x_sx = special_entry_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@220900.4]
  assign package_Anon_io_x_sr = special_entry_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@220900.4]
  assign package_Anon_io_x_pw = special_entry_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@220900.4]
  assign package_Anon_io_x_px = special_entry_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@220900.4]
  assign package_Anon_io_x_pr = special_entry_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@220900.4]
  assign package_Anon_io_x_pal = special_entry_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@220900.4]
  assign package_Anon_io_x_paa = special_entry_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@220900.4]
  assign package_Anon_io_x_eff = special_entry_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@220900.4]
  assign package_Anon_io_x_c = special_entry_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@220900.4]
  assign pmp_io_prv = mpu_priv[1:0]; // @[TLB.scala 193:14:chipyard.TestHarness.RocketConfig.fir@220937.4]
  assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220929.4]
  assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220929.4]
  assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220929.4]
  assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220929.4]
  assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220929.4]
  assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220929.4]
  assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220929.4]
  assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220930.4]
  assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220930.4]
  assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220930.4]
  assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220930.4]
  assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220930.4]
  assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220930.4]
  assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220930.4]
  assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220931.4]
  assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220931.4]
  assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220931.4]
  assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220931.4]
  assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220931.4]
  assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220931.4]
  assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220931.4]
  assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220932.4]
  assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220932.4]
  assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220932.4]
  assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220932.4]
  assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220932.4]
  assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220932.4]
  assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220932.4]
  assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220933.4]
  assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220933.4]
  assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220933.4]
  assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220933.4]
  assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220933.4]
  assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220933.4]
  assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220933.4]
  assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220934.4]
  assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220934.4]
  assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220934.4]
  assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220934.4]
  assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220934.4]
  assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220934.4]
  assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220934.4]
  assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220935.4]
  assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220935.4]
  assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220935.4]
  assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220935.4]
  assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220935.4]
  assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220935.4]
  assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220935.4]
  assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220936.4]
  assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220936.4]
  assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220936.4]
  assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220936.4]
  assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220936.4]
  assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220936.4]
  assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask; // @[TLB.scala 192:14:chipyard.TestHarness.RocketConfig.fir@220936.4]
  assign pmp_io_addr = mpu_physaddr[31:0]; // @[TLB.scala 190:15:chipyard.TestHarness.RocketConfig.fir@220927.4]
  assign package_Anon_1_io_x_ppn = _GEN_35[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221657.4]
  assign package_Anon_1_io_x_u = _GEN_35[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221657.4]
  assign package_Anon_1_io_x_ae = _GEN_35[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221657.4]
  assign package_Anon_1_io_x_sw = _GEN_35[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221657.4]
  assign package_Anon_1_io_x_sx = _GEN_35[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221657.4]
  assign package_Anon_1_io_x_sr = _GEN_35[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221657.4]
  assign package_Anon_1_io_x_pw = _GEN_35[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221657.4]
  assign package_Anon_1_io_x_px = _GEN_35[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221657.4]
  assign package_Anon_1_io_x_pr = _GEN_35[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221657.4]
  assign package_Anon_1_io_x_pal = _GEN_35[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221657.4]
  assign package_Anon_1_io_x_paa = _GEN_35[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221657.4]
  assign package_Anon_1_io_x_eff = _GEN_35[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221657.4]
  assign package_Anon_1_io_x_c = _GEN_35[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221657.4]
  assign package_Anon_2_io_x_ppn = _GEN_39[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221698.4]
  assign package_Anon_2_io_x_u = _GEN_39[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221698.4]
  assign package_Anon_2_io_x_ae = _GEN_39[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221698.4]
  assign package_Anon_2_io_x_sw = _GEN_39[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221698.4]
  assign package_Anon_2_io_x_sx = _GEN_39[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221698.4]
  assign package_Anon_2_io_x_sr = _GEN_39[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221698.4]
  assign package_Anon_2_io_x_pw = _GEN_39[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221698.4]
  assign package_Anon_2_io_x_px = _GEN_39[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221698.4]
  assign package_Anon_2_io_x_pr = _GEN_39[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221698.4]
  assign package_Anon_2_io_x_pal = _GEN_39[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221698.4]
  assign package_Anon_2_io_x_paa = _GEN_39[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221698.4]
  assign package_Anon_2_io_x_eff = _GEN_39[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221698.4]
  assign package_Anon_2_io_x_c = _GEN_39[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221698.4]
  assign package_Anon_3_io_x_ppn = _GEN_43[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221739.4]
  assign package_Anon_3_io_x_u = _GEN_43[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221739.4]
  assign package_Anon_3_io_x_ae = _GEN_43[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221739.4]
  assign package_Anon_3_io_x_sw = _GEN_43[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221739.4]
  assign package_Anon_3_io_x_sx = _GEN_43[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221739.4]
  assign package_Anon_3_io_x_sr = _GEN_43[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221739.4]
  assign package_Anon_3_io_x_pw = _GEN_43[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221739.4]
  assign package_Anon_3_io_x_px = _GEN_43[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221739.4]
  assign package_Anon_3_io_x_pr = _GEN_43[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221739.4]
  assign package_Anon_3_io_x_pal = _GEN_43[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221739.4]
  assign package_Anon_3_io_x_paa = _GEN_43[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221739.4]
  assign package_Anon_3_io_x_eff = _GEN_43[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221739.4]
  assign package_Anon_3_io_x_c = _GEN_43[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221739.4]
  assign package_Anon_4_io_x_ppn = _GEN_47[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221780.4]
  assign package_Anon_4_io_x_u = _GEN_47[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221780.4]
  assign package_Anon_4_io_x_ae = _GEN_47[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221780.4]
  assign package_Anon_4_io_x_sw = _GEN_47[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221780.4]
  assign package_Anon_4_io_x_sx = _GEN_47[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221780.4]
  assign package_Anon_4_io_x_sr = _GEN_47[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221780.4]
  assign package_Anon_4_io_x_pw = _GEN_47[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221780.4]
  assign package_Anon_4_io_x_px = _GEN_47[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221780.4]
  assign package_Anon_4_io_x_pr = _GEN_47[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221780.4]
  assign package_Anon_4_io_x_pal = _GEN_47[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221780.4]
  assign package_Anon_4_io_x_paa = _GEN_47[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221780.4]
  assign package_Anon_4_io_x_eff = _GEN_47[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221780.4]
  assign package_Anon_4_io_x_c = _GEN_47[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221780.4]
  assign package_Anon_5_io_x_ppn = _GEN_51[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221821.4]
  assign package_Anon_5_io_x_u = _GEN_51[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221821.4]
  assign package_Anon_5_io_x_ae = _GEN_51[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221821.4]
  assign package_Anon_5_io_x_sw = _GEN_51[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221821.4]
  assign package_Anon_5_io_x_sx = _GEN_51[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221821.4]
  assign package_Anon_5_io_x_sr = _GEN_51[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221821.4]
  assign package_Anon_5_io_x_pw = _GEN_51[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221821.4]
  assign package_Anon_5_io_x_px = _GEN_51[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221821.4]
  assign package_Anon_5_io_x_pr = _GEN_51[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221821.4]
  assign package_Anon_5_io_x_pal = _GEN_51[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221821.4]
  assign package_Anon_5_io_x_paa = _GEN_51[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221821.4]
  assign package_Anon_5_io_x_eff = _GEN_51[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221821.4]
  assign package_Anon_5_io_x_c = _GEN_51[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221821.4]
  assign package_Anon_6_io_x_ppn = _GEN_55[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221862.4]
  assign package_Anon_6_io_x_u = _GEN_55[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221862.4]
  assign package_Anon_6_io_x_ae = _GEN_55[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221862.4]
  assign package_Anon_6_io_x_sw = _GEN_55[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221862.4]
  assign package_Anon_6_io_x_sx = _GEN_55[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221862.4]
  assign package_Anon_6_io_x_sr = _GEN_55[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221862.4]
  assign package_Anon_6_io_x_pw = _GEN_55[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221862.4]
  assign package_Anon_6_io_x_px = _GEN_55[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221862.4]
  assign package_Anon_6_io_x_pr = _GEN_55[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221862.4]
  assign package_Anon_6_io_x_pal = _GEN_55[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221862.4]
  assign package_Anon_6_io_x_paa = _GEN_55[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221862.4]
  assign package_Anon_6_io_x_eff = _GEN_55[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221862.4]
  assign package_Anon_6_io_x_c = _GEN_55[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221862.4]
  assign package_Anon_7_io_x_ppn = _GEN_59[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221903.4]
  assign package_Anon_7_io_x_u = _GEN_59[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221903.4]
  assign package_Anon_7_io_x_ae = _GEN_59[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221903.4]
  assign package_Anon_7_io_x_sw = _GEN_59[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221903.4]
  assign package_Anon_7_io_x_sx = _GEN_59[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221903.4]
  assign package_Anon_7_io_x_sr = _GEN_59[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221903.4]
  assign package_Anon_7_io_x_pw = _GEN_59[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221903.4]
  assign package_Anon_7_io_x_px = _GEN_59[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221903.4]
  assign package_Anon_7_io_x_pr = _GEN_59[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221903.4]
  assign package_Anon_7_io_x_pal = _GEN_59[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221903.4]
  assign package_Anon_7_io_x_paa = _GEN_59[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221903.4]
  assign package_Anon_7_io_x_eff = _GEN_59[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221903.4]
  assign package_Anon_7_io_x_c = _GEN_59[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221903.4]
  assign package_Anon_8_io_x_ppn = _GEN_63[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221944.4]
  assign package_Anon_8_io_x_u = _GEN_63[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221944.4]
  assign package_Anon_8_io_x_ae = _GEN_63[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221944.4]
  assign package_Anon_8_io_x_sw = _GEN_63[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221944.4]
  assign package_Anon_8_io_x_sx = _GEN_63[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221944.4]
  assign package_Anon_8_io_x_sr = _GEN_63[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221944.4]
  assign package_Anon_8_io_x_pw = _GEN_63[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221944.4]
  assign package_Anon_8_io_x_px = _GEN_63[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221944.4]
  assign package_Anon_8_io_x_pr = _GEN_63[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221944.4]
  assign package_Anon_8_io_x_pal = _GEN_63[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221944.4]
  assign package_Anon_8_io_x_paa = _GEN_63[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221944.4]
  assign package_Anon_8_io_x_eff = _GEN_63[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221944.4]
  assign package_Anon_8_io_x_c = _GEN_63[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221944.4]
  assign package_Anon_9_io_x_ppn = superpage_entries_0_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221984.4]
  assign package_Anon_9_io_x_u = superpage_entries_0_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221984.4]
  assign package_Anon_9_io_x_ae = superpage_entries_0_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221984.4]
  assign package_Anon_9_io_x_sw = superpage_entries_0_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221984.4]
  assign package_Anon_9_io_x_sx = superpage_entries_0_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221984.4]
  assign package_Anon_9_io_x_sr = superpage_entries_0_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221984.4]
  assign package_Anon_9_io_x_pw = superpage_entries_0_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221984.4]
  assign package_Anon_9_io_x_px = superpage_entries_0_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221984.4]
  assign package_Anon_9_io_x_pr = superpage_entries_0_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221984.4]
  assign package_Anon_9_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221984.4]
  assign package_Anon_9_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221984.4]
  assign package_Anon_9_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221984.4]
  assign package_Anon_9_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@221984.4]
  assign package_Anon_10_io_x_ppn = superpage_entries_1_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222037.4]
  assign package_Anon_10_io_x_u = superpage_entries_1_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222037.4]
  assign package_Anon_10_io_x_ae = superpage_entries_1_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222037.4]
  assign package_Anon_10_io_x_sw = superpage_entries_1_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222037.4]
  assign package_Anon_10_io_x_sx = superpage_entries_1_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222037.4]
  assign package_Anon_10_io_x_sr = superpage_entries_1_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222037.4]
  assign package_Anon_10_io_x_pw = superpage_entries_1_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222037.4]
  assign package_Anon_10_io_x_px = superpage_entries_1_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222037.4]
  assign package_Anon_10_io_x_pr = superpage_entries_1_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222037.4]
  assign package_Anon_10_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222037.4]
  assign package_Anon_10_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222037.4]
  assign package_Anon_10_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222037.4]
  assign package_Anon_10_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222037.4]
  assign package_Anon_11_io_x_ppn = superpage_entries_2_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222090.4]
  assign package_Anon_11_io_x_u = superpage_entries_2_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222090.4]
  assign package_Anon_11_io_x_ae = superpage_entries_2_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222090.4]
  assign package_Anon_11_io_x_sw = superpage_entries_2_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222090.4]
  assign package_Anon_11_io_x_sx = superpage_entries_2_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222090.4]
  assign package_Anon_11_io_x_sr = superpage_entries_2_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222090.4]
  assign package_Anon_11_io_x_pw = superpage_entries_2_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222090.4]
  assign package_Anon_11_io_x_px = superpage_entries_2_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222090.4]
  assign package_Anon_11_io_x_pr = superpage_entries_2_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222090.4]
  assign package_Anon_11_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222090.4]
  assign package_Anon_11_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222090.4]
  assign package_Anon_11_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222090.4]
  assign package_Anon_11_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222090.4]
  assign package_Anon_12_io_x_ppn = superpage_entries_3_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222143.4]
  assign package_Anon_12_io_x_u = superpage_entries_3_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222143.4]
  assign package_Anon_12_io_x_ae = superpage_entries_3_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222143.4]
  assign package_Anon_12_io_x_sw = superpage_entries_3_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222143.4]
  assign package_Anon_12_io_x_sx = superpage_entries_3_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222143.4]
  assign package_Anon_12_io_x_sr = superpage_entries_3_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222143.4]
  assign package_Anon_12_io_x_pw = superpage_entries_3_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222143.4]
  assign package_Anon_12_io_x_px = superpage_entries_3_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222143.4]
  assign package_Anon_12_io_x_pr = superpage_entries_3_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222143.4]
  assign package_Anon_12_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222143.4]
  assign package_Anon_12_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222143.4]
  assign package_Anon_12_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222143.4]
  assign package_Anon_12_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222143.4]
  assign package_Anon_13_io_x_ppn = special_entry_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222196.4]
  assign package_Anon_13_io_x_u = special_entry_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222196.4]
  assign package_Anon_13_io_x_ae = special_entry_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222196.4]
  assign package_Anon_13_io_x_sw = special_entry_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222196.4]
  assign package_Anon_13_io_x_sx = special_entry_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222196.4]
  assign package_Anon_13_io_x_sr = special_entry_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222196.4]
  assign package_Anon_13_io_x_pw = special_entry_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222196.4]
  assign package_Anon_13_io_x_px = special_entry_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222196.4]
  assign package_Anon_13_io_x_pr = special_entry_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222196.4]
  assign package_Anon_13_io_x_pal = special_entry_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222196.4]
  assign package_Anon_13_io_x_paa = special_entry_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222196.4]
  assign package_Anon_13_io_x_eff = special_entry_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222196.4]
  assign package_Anon_13_io_x_c = special_entry_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222196.4]
  assign package_Anon_14_io_x_ppn = _GEN_35[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222671.4]
  assign package_Anon_14_io_x_u = _GEN_35[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222671.4]
  assign package_Anon_14_io_x_ae = _GEN_35[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222671.4]
  assign package_Anon_14_io_x_sw = _GEN_35[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222671.4]
  assign package_Anon_14_io_x_sx = _GEN_35[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222671.4]
  assign package_Anon_14_io_x_sr = _GEN_35[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222671.4]
  assign package_Anon_14_io_x_pw = _GEN_35[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222671.4]
  assign package_Anon_14_io_x_px = _GEN_35[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222671.4]
  assign package_Anon_14_io_x_pr = _GEN_35[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222671.4]
  assign package_Anon_14_io_x_pal = _GEN_35[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222671.4]
  assign package_Anon_14_io_x_paa = _GEN_35[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222671.4]
  assign package_Anon_14_io_x_eff = _GEN_35[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222671.4]
  assign package_Anon_14_io_x_c = _GEN_35[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222671.4]
  assign package_Anon_15_io_x_ppn = _GEN_39[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222712.4]
  assign package_Anon_15_io_x_u = _GEN_39[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222712.4]
  assign package_Anon_15_io_x_ae = _GEN_39[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222712.4]
  assign package_Anon_15_io_x_sw = _GEN_39[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222712.4]
  assign package_Anon_15_io_x_sx = _GEN_39[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222712.4]
  assign package_Anon_15_io_x_sr = _GEN_39[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222712.4]
  assign package_Anon_15_io_x_pw = _GEN_39[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222712.4]
  assign package_Anon_15_io_x_px = _GEN_39[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222712.4]
  assign package_Anon_15_io_x_pr = _GEN_39[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222712.4]
  assign package_Anon_15_io_x_pal = _GEN_39[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222712.4]
  assign package_Anon_15_io_x_paa = _GEN_39[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222712.4]
  assign package_Anon_15_io_x_eff = _GEN_39[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222712.4]
  assign package_Anon_15_io_x_c = _GEN_39[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222712.4]
  assign package_Anon_16_io_x_ppn = _GEN_43[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222753.4]
  assign package_Anon_16_io_x_u = _GEN_43[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222753.4]
  assign package_Anon_16_io_x_ae = _GEN_43[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222753.4]
  assign package_Anon_16_io_x_sw = _GEN_43[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222753.4]
  assign package_Anon_16_io_x_sx = _GEN_43[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222753.4]
  assign package_Anon_16_io_x_sr = _GEN_43[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222753.4]
  assign package_Anon_16_io_x_pw = _GEN_43[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222753.4]
  assign package_Anon_16_io_x_px = _GEN_43[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222753.4]
  assign package_Anon_16_io_x_pr = _GEN_43[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222753.4]
  assign package_Anon_16_io_x_pal = _GEN_43[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222753.4]
  assign package_Anon_16_io_x_paa = _GEN_43[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222753.4]
  assign package_Anon_16_io_x_eff = _GEN_43[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222753.4]
  assign package_Anon_16_io_x_c = _GEN_43[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222753.4]
  assign package_Anon_17_io_x_ppn = _GEN_47[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222794.4]
  assign package_Anon_17_io_x_u = _GEN_47[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222794.4]
  assign package_Anon_17_io_x_ae = _GEN_47[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222794.4]
  assign package_Anon_17_io_x_sw = _GEN_47[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222794.4]
  assign package_Anon_17_io_x_sx = _GEN_47[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222794.4]
  assign package_Anon_17_io_x_sr = _GEN_47[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222794.4]
  assign package_Anon_17_io_x_pw = _GEN_47[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222794.4]
  assign package_Anon_17_io_x_px = _GEN_47[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222794.4]
  assign package_Anon_17_io_x_pr = _GEN_47[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222794.4]
  assign package_Anon_17_io_x_pal = _GEN_47[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222794.4]
  assign package_Anon_17_io_x_paa = _GEN_47[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222794.4]
  assign package_Anon_17_io_x_eff = _GEN_47[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222794.4]
  assign package_Anon_17_io_x_c = _GEN_47[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222794.4]
  assign package_Anon_18_io_x_ppn = _GEN_51[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222835.4]
  assign package_Anon_18_io_x_u = _GEN_51[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222835.4]
  assign package_Anon_18_io_x_ae = _GEN_51[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222835.4]
  assign package_Anon_18_io_x_sw = _GEN_51[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222835.4]
  assign package_Anon_18_io_x_sx = _GEN_51[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222835.4]
  assign package_Anon_18_io_x_sr = _GEN_51[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222835.4]
  assign package_Anon_18_io_x_pw = _GEN_51[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222835.4]
  assign package_Anon_18_io_x_px = _GEN_51[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222835.4]
  assign package_Anon_18_io_x_pr = _GEN_51[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222835.4]
  assign package_Anon_18_io_x_pal = _GEN_51[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222835.4]
  assign package_Anon_18_io_x_paa = _GEN_51[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222835.4]
  assign package_Anon_18_io_x_eff = _GEN_51[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222835.4]
  assign package_Anon_18_io_x_c = _GEN_51[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222835.4]
  assign package_Anon_19_io_x_ppn = _GEN_55[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222876.4]
  assign package_Anon_19_io_x_u = _GEN_55[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222876.4]
  assign package_Anon_19_io_x_ae = _GEN_55[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222876.4]
  assign package_Anon_19_io_x_sw = _GEN_55[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222876.4]
  assign package_Anon_19_io_x_sx = _GEN_55[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222876.4]
  assign package_Anon_19_io_x_sr = _GEN_55[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222876.4]
  assign package_Anon_19_io_x_pw = _GEN_55[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222876.4]
  assign package_Anon_19_io_x_px = _GEN_55[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222876.4]
  assign package_Anon_19_io_x_pr = _GEN_55[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222876.4]
  assign package_Anon_19_io_x_pal = _GEN_55[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222876.4]
  assign package_Anon_19_io_x_paa = _GEN_55[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222876.4]
  assign package_Anon_19_io_x_eff = _GEN_55[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222876.4]
  assign package_Anon_19_io_x_c = _GEN_55[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222876.4]
  assign package_Anon_20_io_x_ppn = _GEN_59[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222917.4]
  assign package_Anon_20_io_x_u = _GEN_59[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222917.4]
  assign package_Anon_20_io_x_ae = _GEN_59[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222917.4]
  assign package_Anon_20_io_x_sw = _GEN_59[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222917.4]
  assign package_Anon_20_io_x_sx = _GEN_59[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222917.4]
  assign package_Anon_20_io_x_sr = _GEN_59[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222917.4]
  assign package_Anon_20_io_x_pw = _GEN_59[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222917.4]
  assign package_Anon_20_io_x_px = _GEN_59[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222917.4]
  assign package_Anon_20_io_x_pr = _GEN_59[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222917.4]
  assign package_Anon_20_io_x_pal = _GEN_59[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222917.4]
  assign package_Anon_20_io_x_paa = _GEN_59[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222917.4]
  assign package_Anon_20_io_x_eff = _GEN_59[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222917.4]
  assign package_Anon_20_io_x_c = _GEN_59[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222917.4]
  assign package_Anon_21_io_x_ppn = _GEN_63[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222958.4]
  assign package_Anon_21_io_x_u = _GEN_63[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222958.4]
  assign package_Anon_21_io_x_ae = _GEN_63[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222958.4]
  assign package_Anon_21_io_x_sw = _GEN_63[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222958.4]
  assign package_Anon_21_io_x_sx = _GEN_63[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222958.4]
  assign package_Anon_21_io_x_sr = _GEN_63[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222958.4]
  assign package_Anon_21_io_x_pw = _GEN_63[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222958.4]
  assign package_Anon_21_io_x_px = _GEN_63[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222958.4]
  assign package_Anon_21_io_x_pr = _GEN_63[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222958.4]
  assign package_Anon_21_io_x_pal = _GEN_63[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222958.4]
  assign package_Anon_21_io_x_paa = _GEN_63[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222958.4]
  assign package_Anon_21_io_x_eff = _GEN_63[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222958.4]
  assign package_Anon_21_io_x_c = _GEN_63[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222958.4]
  assign package_Anon_22_io_x_ppn = superpage_entries_0_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222998.4]
  assign package_Anon_22_io_x_u = superpage_entries_0_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222998.4]
  assign package_Anon_22_io_x_ae = superpage_entries_0_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222998.4]
  assign package_Anon_22_io_x_sw = superpage_entries_0_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222998.4]
  assign package_Anon_22_io_x_sx = superpage_entries_0_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222998.4]
  assign package_Anon_22_io_x_sr = superpage_entries_0_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222998.4]
  assign package_Anon_22_io_x_pw = superpage_entries_0_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222998.4]
  assign package_Anon_22_io_x_px = superpage_entries_0_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222998.4]
  assign package_Anon_22_io_x_pr = superpage_entries_0_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222998.4]
  assign package_Anon_22_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222998.4]
  assign package_Anon_22_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222998.4]
  assign package_Anon_22_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222998.4]
  assign package_Anon_22_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@222998.4]
  assign package_Anon_23_io_x_ppn = superpage_entries_1_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223038.4]
  assign package_Anon_23_io_x_u = superpage_entries_1_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223038.4]
  assign package_Anon_23_io_x_ae = superpage_entries_1_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223038.4]
  assign package_Anon_23_io_x_sw = superpage_entries_1_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223038.4]
  assign package_Anon_23_io_x_sx = superpage_entries_1_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223038.4]
  assign package_Anon_23_io_x_sr = superpage_entries_1_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223038.4]
  assign package_Anon_23_io_x_pw = superpage_entries_1_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223038.4]
  assign package_Anon_23_io_x_px = superpage_entries_1_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223038.4]
  assign package_Anon_23_io_x_pr = superpage_entries_1_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223038.4]
  assign package_Anon_23_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223038.4]
  assign package_Anon_23_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223038.4]
  assign package_Anon_23_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223038.4]
  assign package_Anon_23_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223038.4]
  assign package_Anon_24_io_x_ppn = superpage_entries_2_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223078.4]
  assign package_Anon_24_io_x_u = superpage_entries_2_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223078.4]
  assign package_Anon_24_io_x_ae = superpage_entries_2_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223078.4]
  assign package_Anon_24_io_x_sw = superpage_entries_2_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223078.4]
  assign package_Anon_24_io_x_sx = superpage_entries_2_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223078.4]
  assign package_Anon_24_io_x_sr = superpage_entries_2_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223078.4]
  assign package_Anon_24_io_x_pw = superpage_entries_2_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223078.4]
  assign package_Anon_24_io_x_px = superpage_entries_2_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223078.4]
  assign package_Anon_24_io_x_pr = superpage_entries_2_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223078.4]
  assign package_Anon_24_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223078.4]
  assign package_Anon_24_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223078.4]
  assign package_Anon_24_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223078.4]
  assign package_Anon_24_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223078.4]
  assign package_Anon_25_io_x_ppn = superpage_entries_3_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223118.4]
  assign package_Anon_25_io_x_u = superpage_entries_3_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223118.4]
  assign package_Anon_25_io_x_ae = superpage_entries_3_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223118.4]
  assign package_Anon_25_io_x_sw = superpage_entries_3_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223118.4]
  assign package_Anon_25_io_x_sx = superpage_entries_3_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223118.4]
  assign package_Anon_25_io_x_sr = superpage_entries_3_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223118.4]
  assign package_Anon_25_io_x_pw = superpage_entries_3_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223118.4]
  assign package_Anon_25_io_x_px = superpage_entries_3_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223118.4]
  assign package_Anon_25_io_x_pr = superpage_entries_3_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223118.4]
  assign package_Anon_25_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223118.4]
  assign package_Anon_25_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223118.4]
  assign package_Anon_25_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223118.4]
  assign package_Anon_25_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223118.4]
  assign package_Anon_26_io_x_ppn = special_entry_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223158.4]
  assign package_Anon_26_io_x_u = special_entry_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223158.4]
  assign package_Anon_26_io_x_ae = special_entry_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223158.4]
  assign package_Anon_26_io_x_sw = special_entry_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223158.4]
  assign package_Anon_26_io_x_sx = special_entry_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223158.4]
  assign package_Anon_26_io_x_sr = special_entry_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223158.4]
  assign package_Anon_26_io_x_pw = special_entry_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223158.4]
  assign package_Anon_26_io_x_px = special_entry_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223158.4]
  assign package_Anon_26_io_x_pr = special_entry_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223158.4]
  assign package_Anon_26_io_x_pal = special_entry_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223158.4]
  assign package_Anon_26_io_x_paa = special_entry_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223158.4]
  assign package_Anon_26_io_x_eff = special_entry_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223158.4]
  assign package_Anon_26_io_x_c = special_entry_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223158.4]
  assign package_Anon_27_io_x_ppn = _GEN_35[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223199.4]
  assign package_Anon_27_io_x_u = _GEN_35[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223199.4]
  assign package_Anon_27_io_x_ae = _GEN_35[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223199.4]
  assign package_Anon_27_io_x_sw = _GEN_35[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223199.4]
  assign package_Anon_27_io_x_sx = _GEN_35[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223199.4]
  assign package_Anon_27_io_x_sr = _GEN_35[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223199.4]
  assign package_Anon_27_io_x_pw = _GEN_35[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223199.4]
  assign package_Anon_27_io_x_px = _GEN_35[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223199.4]
  assign package_Anon_27_io_x_pr = _GEN_35[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223199.4]
  assign package_Anon_27_io_x_pal = _GEN_35[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223199.4]
  assign package_Anon_27_io_x_paa = _GEN_35[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223199.4]
  assign package_Anon_27_io_x_eff = _GEN_35[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223199.4]
  assign package_Anon_27_io_x_c = _GEN_35[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223199.4]
  assign package_Anon_28_io_x_ppn = _GEN_39[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223240.4]
  assign package_Anon_28_io_x_u = _GEN_39[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223240.4]
  assign package_Anon_28_io_x_ae = _GEN_39[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223240.4]
  assign package_Anon_28_io_x_sw = _GEN_39[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223240.4]
  assign package_Anon_28_io_x_sx = _GEN_39[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223240.4]
  assign package_Anon_28_io_x_sr = _GEN_39[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223240.4]
  assign package_Anon_28_io_x_pw = _GEN_39[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223240.4]
  assign package_Anon_28_io_x_px = _GEN_39[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223240.4]
  assign package_Anon_28_io_x_pr = _GEN_39[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223240.4]
  assign package_Anon_28_io_x_pal = _GEN_39[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223240.4]
  assign package_Anon_28_io_x_paa = _GEN_39[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223240.4]
  assign package_Anon_28_io_x_eff = _GEN_39[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223240.4]
  assign package_Anon_28_io_x_c = _GEN_39[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223240.4]
  assign package_Anon_29_io_x_ppn = _GEN_43[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223281.4]
  assign package_Anon_29_io_x_u = _GEN_43[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223281.4]
  assign package_Anon_29_io_x_ae = _GEN_43[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223281.4]
  assign package_Anon_29_io_x_sw = _GEN_43[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223281.4]
  assign package_Anon_29_io_x_sx = _GEN_43[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223281.4]
  assign package_Anon_29_io_x_sr = _GEN_43[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223281.4]
  assign package_Anon_29_io_x_pw = _GEN_43[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223281.4]
  assign package_Anon_29_io_x_px = _GEN_43[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223281.4]
  assign package_Anon_29_io_x_pr = _GEN_43[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223281.4]
  assign package_Anon_29_io_x_pal = _GEN_43[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223281.4]
  assign package_Anon_29_io_x_paa = _GEN_43[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223281.4]
  assign package_Anon_29_io_x_eff = _GEN_43[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223281.4]
  assign package_Anon_29_io_x_c = _GEN_43[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223281.4]
  assign package_Anon_30_io_x_ppn = _GEN_47[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223322.4]
  assign package_Anon_30_io_x_u = _GEN_47[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223322.4]
  assign package_Anon_30_io_x_ae = _GEN_47[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223322.4]
  assign package_Anon_30_io_x_sw = _GEN_47[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223322.4]
  assign package_Anon_30_io_x_sx = _GEN_47[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223322.4]
  assign package_Anon_30_io_x_sr = _GEN_47[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223322.4]
  assign package_Anon_30_io_x_pw = _GEN_47[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223322.4]
  assign package_Anon_30_io_x_px = _GEN_47[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223322.4]
  assign package_Anon_30_io_x_pr = _GEN_47[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223322.4]
  assign package_Anon_30_io_x_pal = _GEN_47[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223322.4]
  assign package_Anon_30_io_x_paa = _GEN_47[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223322.4]
  assign package_Anon_30_io_x_eff = _GEN_47[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223322.4]
  assign package_Anon_30_io_x_c = _GEN_47[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223322.4]
  assign package_Anon_31_io_x_ppn = _GEN_51[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223363.4]
  assign package_Anon_31_io_x_u = _GEN_51[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223363.4]
  assign package_Anon_31_io_x_ae = _GEN_51[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223363.4]
  assign package_Anon_31_io_x_sw = _GEN_51[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223363.4]
  assign package_Anon_31_io_x_sx = _GEN_51[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223363.4]
  assign package_Anon_31_io_x_sr = _GEN_51[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223363.4]
  assign package_Anon_31_io_x_pw = _GEN_51[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223363.4]
  assign package_Anon_31_io_x_px = _GEN_51[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223363.4]
  assign package_Anon_31_io_x_pr = _GEN_51[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223363.4]
  assign package_Anon_31_io_x_pal = _GEN_51[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223363.4]
  assign package_Anon_31_io_x_paa = _GEN_51[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223363.4]
  assign package_Anon_31_io_x_eff = _GEN_51[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223363.4]
  assign package_Anon_31_io_x_c = _GEN_51[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223363.4]
  assign package_Anon_32_io_x_ppn = _GEN_55[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223404.4]
  assign package_Anon_32_io_x_u = _GEN_55[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223404.4]
  assign package_Anon_32_io_x_ae = _GEN_55[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223404.4]
  assign package_Anon_32_io_x_sw = _GEN_55[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223404.4]
  assign package_Anon_32_io_x_sx = _GEN_55[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223404.4]
  assign package_Anon_32_io_x_sr = _GEN_55[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223404.4]
  assign package_Anon_32_io_x_pw = _GEN_55[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223404.4]
  assign package_Anon_32_io_x_px = _GEN_55[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223404.4]
  assign package_Anon_32_io_x_pr = _GEN_55[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223404.4]
  assign package_Anon_32_io_x_pal = _GEN_55[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223404.4]
  assign package_Anon_32_io_x_paa = _GEN_55[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223404.4]
  assign package_Anon_32_io_x_eff = _GEN_55[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223404.4]
  assign package_Anon_32_io_x_c = _GEN_55[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223404.4]
  assign package_Anon_33_io_x_ppn = _GEN_59[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223445.4]
  assign package_Anon_33_io_x_u = _GEN_59[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223445.4]
  assign package_Anon_33_io_x_ae = _GEN_59[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223445.4]
  assign package_Anon_33_io_x_sw = _GEN_59[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223445.4]
  assign package_Anon_33_io_x_sx = _GEN_59[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223445.4]
  assign package_Anon_33_io_x_sr = _GEN_59[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223445.4]
  assign package_Anon_33_io_x_pw = _GEN_59[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223445.4]
  assign package_Anon_33_io_x_px = _GEN_59[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223445.4]
  assign package_Anon_33_io_x_pr = _GEN_59[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223445.4]
  assign package_Anon_33_io_x_pal = _GEN_59[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223445.4]
  assign package_Anon_33_io_x_paa = _GEN_59[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223445.4]
  assign package_Anon_33_io_x_eff = _GEN_59[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223445.4]
  assign package_Anon_33_io_x_c = _GEN_59[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223445.4]
  assign package_Anon_34_io_x_ppn = _GEN_63[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223486.4]
  assign package_Anon_34_io_x_u = _GEN_63[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223486.4]
  assign package_Anon_34_io_x_ae = _GEN_63[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223486.4]
  assign package_Anon_34_io_x_sw = _GEN_63[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223486.4]
  assign package_Anon_34_io_x_sx = _GEN_63[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223486.4]
  assign package_Anon_34_io_x_sr = _GEN_63[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223486.4]
  assign package_Anon_34_io_x_pw = _GEN_63[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223486.4]
  assign package_Anon_34_io_x_px = _GEN_63[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223486.4]
  assign package_Anon_34_io_x_pr = _GEN_63[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223486.4]
  assign package_Anon_34_io_x_pal = _GEN_63[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223486.4]
  assign package_Anon_34_io_x_paa = _GEN_63[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223486.4]
  assign package_Anon_34_io_x_eff = _GEN_63[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223486.4]
  assign package_Anon_34_io_x_c = _GEN_63[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223486.4]
  assign package_Anon_35_io_x_ppn = superpage_entries_0_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223526.4]
  assign package_Anon_35_io_x_u = superpage_entries_0_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223526.4]
  assign package_Anon_35_io_x_ae = superpage_entries_0_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223526.4]
  assign package_Anon_35_io_x_sw = superpage_entries_0_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223526.4]
  assign package_Anon_35_io_x_sx = superpage_entries_0_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223526.4]
  assign package_Anon_35_io_x_sr = superpage_entries_0_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223526.4]
  assign package_Anon_35_io_x_pw = superpage_entries_0_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223526.4]
  assign package_Anon_35_io_x_px = superpage_entries_0_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223526.4]
  assign package_Anon_35_io_x_pr = superpage_entries_0_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223526.4]
  assign package_Anon_35_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223526.4]
  assign package_Anon_35_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223526.4]
  assign package_Anon_35_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223526.4]
  assign package_Anon_35_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223526.4]
  assign package_Anon_36_io_x_ppn = superpage_entries_1_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223566.4]
  assign package_Anon_36_io_x_u = superpage_entries_1_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223566.4]
  assign package_Anon_36_io_x_ae = superpage_entries_1_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223566.4]
  assign package_Anon_36_io_x_sw = superpage_entries_1_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223566.4]
  assign package_Anon_36_io_x_sx = superpage_entries_1_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223566.4]
  assign package_Anon_36_io_x_sr = superpage_entries_1_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223566.4]
  assign package_Anon_36_io_x_pw = superpage_entries_1_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223566.4]
  assign package_Anon_36_io_x_px = superpage_entries_1_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223566.4]
  assign package_Anon_36_io_x_pr = superpage_entries_1_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223566.4]
  assign package_Anon_36_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223566.4]
  assign package_Anon_36_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223566.4]
  assign package_Anon_36_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223566.4]
  assign package_Anon_36_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223566.4]
  assign package_Anon_37_io_x_ppn = superpage_entries_2_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223606.4]
  assign package_Anon_37_io_x_u = superpage_entries_2_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223606.4]
  assign package_Anon_37_io_x_ae = superpage_entries_2_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223606.4]
  assign package_Anon_37_io_x_sw = superpage_entries_2_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223606.4]
  assign package_Anon_37_io_x_sx = superpage_entries_2_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223606.4]
  assign package_Anon_37_io_x_sr = superpage_entries_2_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223606.4]
  assign package_Anon_37_io_x_pw = superpage_entries_2_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223606.4]
  assign package_Anon_37_io_x_px = superpage_entries_2_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223606.4]
  assign package_Anon_37_io_x_pr = superpage_entries_2_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223606.4]
  assign package_Anon_37_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223606.4]
  assign package_Anon_37_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223606.4]
  assign package_Anon_37_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223606.4]
  assign package_Anon_37_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223606.4]
  assign package_Anon_38_io_x_ppn = superpage_entries_3_data_0[33:14]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223646.4]
  assign package_Anon_38_io_x_u = superpage_entries_3_data_0[13]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223646.4]
  assign package_Anon_38_io_x_ae = superpage_entries_3_data_0[11]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223646.4]
  assign package_Anon_38_io_x_sw = superpage_entries_3_data_0[10]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223646.4]
  assign package_Anon_38_io_x_sx = superpage_entries_3_data_0[9]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223646.4]
  assign package_Anon_38_io_x_sr = superpage_entries_3_data_0[8]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223646.4]
  assign package_Anon_38_io_x_pw = superpage_entries_3_data_0[7]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223646.4]
  assign package_Anon_38_io_x_px = superpage_entries_3_data_0[6]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223646.4]
  assign package_Anon_38_io_x_pr = superpage_entries_3_data_0[5]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223646.4]
  assign package_Anon_38_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223646.4]
  assign package_Anon_38_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223646.4]
  assign package_Anon_38_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223646.4]
  assign package_Anon_38_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 220:14:chipyard.TestHarness.RocketConfig.fir@223646.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_tag = _RAND_0[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_data_0 = _RAND_1[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_data_1 = _RAND_2[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_data_2 = _RAND_3[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_data_3 = _RAND_4[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_valid_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_valid_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_valid_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_valid_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_1_tag = _RAND_9[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_1_data_0 = _RAND_10[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_1_data_1 = _RAND_11[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_1_data_2 = _RAND_12[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_1_data_3 = _RAND_13[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_1_valid_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_1_valid_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_1_valid_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_1_valid_3 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sectored_entries_2_tag = _RAND_18[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  sectored_entries_2_data_0 = _RAND_19[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  sectored_entries_2_data_1 = _RAND_20[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  sectored_entries_2_data_2 = _RAND_21[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  sectored_entries_2_data_3 = _RAND_22[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sectored_entries_2_valid_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sectored_entries_2_valid_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sectored_entries_2_valid_2 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sectored_entries_2_valid_3 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sectored_entries_3_tag = _RAND_27[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  sectored_entries_3_data_0 = _RAND_28[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  sectored_entries_3_data_1 = _RAND_29[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  sectored_entries_3_data_2 = _RAND_30[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  sectored_entries_3_data_3 = _RAND_31[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  sectored_entries_3_valid_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  sectored_entries_3_valid_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  sectored_entries_3_valid_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  sectored_entries_3_valid_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  sectored_entries_4_tag = _RAND_36[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  sectored_entries_4_data_0 = _RAND_37[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  sectored_entries_4_data_1 = _RAND_38[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  sectored_entries_4_data_2 = _RAND_39[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  sectored_entries_4_data_3 = _RAND_40[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  sectored_entries_4_valid_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  sectored_entries_4_valid_1 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  sectored_entries_4_valid_2 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  sectored_entries_4_valid_3 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  sectored_entries_5_tag = _RAND_45[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  sectored_entries_5_data_0 = _RAND_46[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  sectored_entries_5_data_1 = _RAND_47[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  sectored_entries_5_data_2 = _RAND_48[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  sectored_entries_5_data_3 = _RAND_49[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  sectored_entries_5_valid_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  sectored_entries_5_valid_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  sectored_entries_5_valid_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  sectored_entries_5_valid_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  sectored_entries_6_tag = _RAND_54[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  sectored_entries_6_data_0 = _RAND_55[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {2{`RANDOM}};
  sectored_entries_6_data_1 = _RAND_56[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  sectored_entries_6_data_2 = _RAND_57[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  sectored_entries_6_data_3 = _RAND_58[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  sectored_entries_6_valid_0 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  sectored_entries_6_valid_1 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  sectored_entries_6_valid_2 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  sectored_entries_6_valid_3 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  sectored_entries_7_tag = _RAND_63[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {2{`RANDOM}};
  sectored_entries_7_data_0 = _RAND_64[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  sectored_entries_7_data_1 = _RAND_65[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  sectored_entries_7_data_2 = _RAND_66[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  sectored_entries_7_data_3 = _RAND_67[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  sectored_entries_7_valid_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  sectored_entries_7_valid_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  sectored_entries_7_valid_2 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  sectored_entries_7_valid_3 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  superpage_entries_0_level = _RAND_72[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  superpage_entries_0_tag = _RAND_73[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_74[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  superpage_entries_1_level = _RAND_76[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  superpage_entries_1_tag = _RAND_77[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_78[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  superpage_entries_2_level = _RAND_80[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  superpage_entries_2_tag = _RAND_81[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{`RANDOM}};
  superpage_entries_2_data_0 = _RAND_82[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  superpage_entries_2_valid_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  superpage_entries_3_level = _RAND_84[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  superpage_entries_3_tag = _RAND_85[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{`RANDOM}};
  superpage_entries_3_data_0 = _RAND_86[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  superpage_entries_3_valid_0 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  special_entry_level = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  special_entry_tag = _RAND_89[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_90[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  state = _RAND_92[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  r_refill_tag = _RAND_93[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_94[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_95[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  r_sectored_hit_addr = _RAND_96[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  r_sectored_hit = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_2015 = _RAND_98[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_2016 = _RAND_99[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1098) begin
            sectored_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1098) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_0 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1098) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_1 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1098) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_2 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1098) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_0_data_3 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_3735) begin
      sectored_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2369) begin
          if (sectored_entries_0_data_0[0]) begin
            sectored_entries_0_valid_0 <= 1'h0;
          end else if (_T_389) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_0_valid_0 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1098) begin
                    sectored_entries_0_valid_0 <= _GEN_84;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1098) begin
                  sectored_entries_0_valid_0 <= _GEN_84;
                end
              end
            end
          end
        end else if (_T_389) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_0_valid_0 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1098) begin
                  sectored_entries_0_valid_0 <= _GEN_84;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1098) begin
                sectored_entries_0_valid_0 <= _GEN_84;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_0 <= _GEN_652;
      end
    end else begin
      sectored_entries_0_valid_0 <= _GEN_472;
    end
    if (_T_3735) begin
      sectored_entries_0_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2369) begin
          if (sectored_entries_0_data_1[0]) begin
            sectored_entries_0_valid_1 <= 1'h0;
          end else if (_T_389) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_0_valid_1 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1098) begin
                    sectored_entries_0_valid_1 <= _GEN_85;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1098) begin
                  sectored_entries_0_valid_1 <= _GEN_85;
                end
              end
            end
          end
        end else if (_T_389) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_0_valid_1 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1098) begin
                  sectored_entries_0_valid_1 <= _GEN_85;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1098) begin
                sectored_entries_0_valid_1 <= _GEN_85;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_1 <= _GEN_653;
      end
    end else begin
      sectored_entries_0_valid_1 <= _GEN_473;
    end
    if (_T_3735) begin
      sectored_entries_0_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2369) begin
          if (sectored_entries_0_data_2[0]) begin
            sectored_entries_0_valid_2 <= 1'h0;
          end else if (_T_389) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_0_valid_2 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1098) begin
                    sectored_entries_0_valid_2 <= _GEN_86;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1098) begin
                  sectored_entries_0_valid_2 <= _GEN_86;
                end
              end
            end
          end
        end else if (_T_389) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_0_valid_2 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1098) begin
                  sectored_entries_0_valid_2 <= _GEN_86;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1098) begin
                sectored_entries_0_valid_2 <= _GEN_86;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_2 <= _GEN_654;
      end
    end else begin
      sectored_entries_0_valid_2 <= _GEN_474;
    end
    if (_T_3735) begin
      sectored_entries_0_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2369) begin
          if (sectored_entries_0_data_3[0]) begin
            sectored_entries_0_valid_3 <= 1'h0;
          end else if (_T_389) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_0_valid_3 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1098) begin
                    sectored_entries_0_valid_3 <= _GEN_87;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1098) begin
                  sectored_entries_0_valid_3 <= _GEN_87;
                end
              end
            end
          end
        end else if (_T_389) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_0_valid_3 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1098) begin
                  sectored_entries_0_valid_3 <= _GEN_87;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1098) begin
                sectored_entries_0_valid_3 <= _GEN_87;
              end
            end
          end
        end
      end else begin
        sectored_entries_0_valid_3 <= _GEN_655;
      end
    end else begin
      sectored_entries_0_valid_3 <= _GEN_475;
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1115) begin
            sectored_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1115) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_0 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1115) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_1 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1115) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_2 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1115) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_1_data_3 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_3735) begin
      sectored_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2516) begin
          if (sectored_entries_1_data_0[0]) begin
            sectored_entries_1_valid_0 <= 1'h0;
          end else if (_T_395) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_1_valid_0 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1115) begin
                    sectored_entries_1_valid_0 <= _GEN_106;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1115) begin
                  sectored_entries_1_valid_0 <= _GEN_106;
                end
              end
            end
          end
        end else if (_T_395) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_1_valid_0 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1115) begin
                  sectored_entries_1_valid_0 <= _GEN_106;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1115) begin
                sectored_entries_1_valid_0 <= _GEN_106;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_0 <= _GEN_680;
      end
    end else begin
      sectored_entries_1_valid_0 <= _GEN_482;
    end
    if (_T_3735) begin
      sectored_entries_1_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2516) begin
          if (sectored_entries_1_data_1[0]) begin
            sectored_entries_1_valid_1 <= 1'h0;
          end else if (_T_395) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_1_valid_1 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1115) begin
                    sectored_entries_1_valid_1 <= _GEN_107;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1115) begin
                  sectored_entries_1_valid_1 <= _GEN_107;
                end
              end
            end
          end
        end else if (_T_395) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_1_valid_1 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1115) begin
                  sectored_entries_1_valid_1 <= _GEN_107;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1115) begin
                sectored_entries_1_valid_1 <= _GEN_107;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_1 <= _GEN_681;
      end
    end else begin
      sectored_entries_1_valid_1 <= _GEN_483;
    end
    if (_T_3735) begin
      sectored_entries_1_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2516) begin
          if (sectored_entries_1_data_2[0]) begin
            sectored_entries_1_valid_2 <= 1'h0;
          end else if (_T_395) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_1_valid_2 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1115) begin
                    sectored_entries_1_valid_2 <= _GEN_108;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1115) begin
                  sectored_entries_1_valid_2 <= _GEN_108;
                end
              end
            end
          end
        end else if (_T_395) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_1_valid_2 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1115) begin
                  sectored_entries_1_valid_2 <= _GEN_108;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1115) begin
                sectored_entries_1_valid_2 <= _GEN_108;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_2 <= _GEN_682;
      end
    end else begin
      sectored_entries_1_valid_2 <= _GEN_484;
    end
    if (_T_3735) begin
      sectored_entries_1_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2516) begin
          if (sectored_entries_1_data_3[0]) begin
            sectored_entries_1_valid_3 <= 1'h0;
          end else if (_T_395) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_1_valid_3 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1115) begin
                    sectored_entries_1_valid_3 <= _GEN_109;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1115) begin
                  sectored_entries_1_valid_3 <= _GEN_109;
                end
              end
            end
          end
        end else if (_T_395) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_1_valid_3 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1115) begin
                  sectored_entries_1_valid_3 <= _GEN_109;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1115) begin
                sectored_entries_1_valid_3 <= _GEN_109;
              end
            end
          end
        end
      end else begin
        sectored_entries_1_valid_3 <= _GEN_683;
      end
    end else begin
      sectored_entries_1_valid_3 <= _GEN_485;
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1132) begin
            sectored_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1132) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_0 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1132) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_1 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1132) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_2 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1132) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_2_data_3 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_3735) begin
      sectored_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2663) begin
          if (sectored_entries_2_data_0[0]) begin
            sectored_entries_2_valid_0 <= 1'h0;
          end else if (_T_401) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_2_valid_0 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1132) begin
                    sectored_entries_2_valid_0 <= _GEN_128;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1132) begin
                  sectored_entries_2_valid_0 <= _GEN_128;
                end
              end
            end
          end
        end else if (_T_401) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_2_valid_0 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1132) begin
                  sectored_entries_2_valid_0 <= _GEN_128;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1132) begin
                sectored_entries_2_valid_0 <= _GEN_128;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_0 <= _GEN_708;
      end
    end else begin
      sectored_entries_2_valid_0 <= _GEN_492;
    end
    if (_T_3735) begin
      sectored_entries_2_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2663) begin
          if (sectored_entries_2_data_1[0]) begin
            sectored_entries_2_valid_1 <= 1'h0;
          end else if (_T_401) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_2_valid_1 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1132) begin
                    sectored_entries_2_valid_1 <= _GEN_129;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1132) begin
                  sectored_entries_2_valid_1 <= _GEN_129;
                end
              end
            end
          end
        end else if (_T_401) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_2_valid_1 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1132) begin
                  sectored_entries_2_valid_1 <= _GEN_129;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1132) begin
                sectored_entries_2_valid_1 <= _GEN_129;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_1 <= _GEN_709;
      end
    end else begin
      sectored_entries_2_valid_1 <= _GEN_493;
    end
    if (_T_3735) begin
      sectored_entries_2_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2663) begin
          if (sectored_entries_2_data_2[0]) begin
            sectored_entries_2_valid_2 <= 1'h0;
          end else if (_T_401) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_2_valid_2 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1132) begin
                    sectored_entries_2_valid_2 <= _GEN_130;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1132) begin
                  sectored_entries_2_valid_2 <= _GEN_130;
                end
              end
            end
          end
        end else if (_T_401) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_2_valid_2 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1132) begin
                  sectored_entries_2_valid_2 <= _GEN_130;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1132) begin
                sectored_entries_2_valid_2 <= _GEN_130;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_2 <= _GEN_710;
      end
    end else begin
      sectored_entries_2_valid_2 <= _GEN_494;
    end
    if (_T_3735) begin
      sectored_entries_2_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2663) begin
          if (sectored_entries_2_data_3[0]) begin
            sectored_entries_2_valid_3 <= 1'h0;
          end else if (_T_401) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_2_valid_3 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1132) begin
                    sectored_entries_2_valid_3 <= _GEN_131;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1132) begin
                  sectored_entries_2_valid_3 <= _GEN_131;
                end
              end
            end
          end
        end else if (_T_401) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_2_valid_3 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1132) begin
                  sectored_entries_2_valid_3 <= _GEN_131;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1132) begin
                sectored_entries_2_valid_3 <= _GEN_131;
              end
            end
          end
        end
      end else begin
        sectored_entries_2_valid_3 <= _GEN_711;
      end
    end else begin
      sectored_entries_2_valid_3 <= _GEN_495;
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1149) begin
            sectored_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1149) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_0 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1149) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_1 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1149) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_2 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1149) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_3_data_3 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_3735) begin
      sectored_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2810) begin
          if (sectored_entries_3_data_0[0]) begin
            sectored_entries_3_valid_0 <= 1'h0;
          end else if (_T_407) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_3_valid_0 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1149) begin
                    sectored_entries_3_valid_0 <= _GEN_150;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1149) begin
                  sectored_entries_3_valid_0 <= _GEN_150;
                end
              end
            end
          end
        end else if (_T_407) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_3_valid_0 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1149) begin
                  sectored_entries_3_valid_0 <= _GEN_150;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1149) begin
                sectored_entries_3_valid_0 <= _GEN_150;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_0 <= _GEN_736;
      end
    end else begin
      sectored_entries_3_valid_0 <= _GEN_502;
    end
    if (_T_3735) begin
      sectored_entries_3_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2810) begin
          if (sectored_entries_3_data_1[0]) begin
            sectored_entries_3_valid_1 <= 1'h0;
          end else if (_T_407) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_3_valid_1 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1149) begin
                    sectored_entries_3_valid_1 <= _GEN_151;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1149) begin
                  sectored_entries_3_valid_1 <= _GEN_151;
                end
              end
            end
          end
        end else if (_T_407) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_3_valid_1 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1149) begin
                  sectored_entries_3_valid_1 <= _GEN_151;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1149) begin
                sectored_entries_3_valid_1 <= _GEN_151;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_1 <= _GEN_737;
      end
    end else begin
      sectored_entries_3_valid_1 <= _GEN_503;
    end
    if (_T_3735) begin
      sectored_entries_3_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2810) begin
          if (sectored_entries_3_data_2[0]) begin
            sectored_entries_3_valid_2 <= 1'h0;
          end else if (_T_407) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_3_valid_2 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1149) begin
                    sectored_entries_3_valid_2 <= _GEN_152;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1149) begin
                  sectored_entries_3_valid_2 <= _GEN_152;
                end
              end
            end
          end
        end else if (_T_407) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_3_valid_2 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1149) begin
                  sectored_entries_3_valid_2 <= _GEN_152;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1149) begin
                sectored_entries_3_valid_2 <= _GEN_152;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_2 <= _GEN_738;
      end
    end else begin
      sectored_entries_3_valid_2 <= _GEN_504;
    end
    if (_T_3735) begin
      sectored_entries_3_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2810) begin
          if (sectored_entries_3_data_3[0]) begin
            sectored_entries_3_valid_3 <= 1'h0;
          end else if (_T_407) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_3_valid_3 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1149) begin
                    sectored_entries_3_valid_3 <= _GEN_153;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1149) begin
                  sectored_entries_3_valid_3 <= _GEN_153;
                end
              end
            end
          end
        end else if (_T_407) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_3_valid_3 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1149) begin
                  sectored_entries_3_valid_3 <= _GEN_153;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1149) begin
                sectored_entries_3_valid_3 <= _GEN_153;
              end
            end
          end
        end
      end else begin
        sectored_entries_3_valid_3 <= _GEN_739;
      end
    end else begin
      sectored_entries_3_valid_3 <= _GEN_505;
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1166) begin
            sectored_entries_4_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1166) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_0 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1166) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_1 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1166) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_2 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1166) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_4_data_3 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_3735) begin
      sectored_entries_4_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2957) begin
          if (sectored_entries_4_data_0[0]) begin
            sectored_entries_4_valid_0 <= 1'h0;
          end else if (_T_413) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_4_valid_0 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1166) begin
                    sectored_entries_4_valid_0 <= _GEN_172;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1166) begin
                  sectored_entries_4_valid_0 <= _GEN_172;
                end
              end
            end
          end
        end else if (_T_413) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_4_valid_0 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1166) begin
                  sectored_entries_4_valid_0 <= _GEN_172;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1166) begin
                sectored_entries_4_valid_0 <= _GEN_172;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_0 <= _GEN_764;
      end
    end else begin
      sectored_entries_4_valid_0 <= _GEN_512;
    end
    if (_T_3735) begin
      sectored_entries_4_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2957) begin
          if (sectored_entries_4_data_1[0]) begin
            sectored_entries_4_valid_1 <= 1'h0;
          end else if (_T_413) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_4_valid_1 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1166) begin
                    sectored_entries_4_valid_1 <= _GEN_173;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1166) begin
                  sectored_entries_4_valid_1 <= _GEN_173;
                end
              end
            end
          end
        end else if (_T_413) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_4_valid_1 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1166) begin
                  sectored_entries_4_valid_1 <= _GEN_173;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1166) begin
                sectored_entries_4_valid_1 <= _GEN_173;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_1 <= _GEN_765;
      end
    end else begin
      sectored_entries_4_valid_1 <= _GEN_513;
    end
    if (_T_3735) begin
      sectored_entries_4_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2957) begin
          if (sectored_entries_4_data_2[0]) begin
            sectored_entries_4_valid_2 <= 1'h0;
          end else if (_T_413) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_4_valid_2 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1166) begin
                    sectored_entries_4_valid_2 <= _GEN_174;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1166) begin
                  sectored_entries_4_valid_2 <= _GEN_174;
                end
              end
            end
          end
        end else if (_T_413) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_4_valid_2 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1166) begin
                  sectored_entries_4_valid_2 <= _GEN_174;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1166) begin
                sectored_entries_4_valid_2 <= _GEN_174;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_2 <= _GEN_766;
      end
    end else begin
      sectored_entries_4_valid_2 <= _GEN_514;
    end
    if (_T_3735) begin
      sectored_entries_4_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_2957) begin
          if (sectored_entries_4_data_3[0]) begin
            sectored_entries_4_valid_3 <= 1'h0;
          end else if (_T_413) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_4_valid_3 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1166) begin
                    sectored_entries_4_valid_3 <= _GEN_175;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1166) begin
                  sectored_entries_4_valid_3 <= _GEN_175;
                end
              end
            end
          end
        end else if (_T_413) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_4_valid_3 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1166) begin
                  sectored_entries_4_valid_3 <= _GEN_175;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1166) begin
                sectored_entries_4_valid_3 <= _GEN_175;
              end
            end
          end
        end
      end else begin
        sectored_entries_4_valid_3 <= _GEN_767;
      end
    end else begin
      sectored_entries_4_valid_3 <= _GEN_515;
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1183) begin
            sectored_entries_5_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1183) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_0 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1183) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_1 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1183) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_2 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1183) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_5_data_3 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_3735) begin
      sectored_entries_5_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3104) begin
          if (sectored_entries_5_data_0[0]) begin
            sectored_entries_5_valid_0 <= 1'h0;
          end else if (_T_419) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_5_valid_0 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1183) begin
                    sectored_entries_5_valid_0 <= _GEN_194;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1183) begin
                  sectored_entries_5_valid_0 <= _GEN_194;
                end
              end
            end
          end
        end else if (_T_419) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_5_valid_0 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1183) begin
                  sectored_entries_5_valid_0 <= _GEN_194;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1183) begin
                sectored_entries_5_valid_0 <= _GEN_194;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_0 <= _GEN_792;
      end
    end else begin
      sectored_entries_5_valid_0 <= _GEN_522;
    end
    if (_T_3735) begin
      sectored_entries_5_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3104) begin
          if (sectored_entries_5_data_1[0]) begin
            sectored_entries_5_valid_1 <= 1'h0;
          end else if (_T_419) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_5_valid_1 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1183) begin
                    sectored_entries_5_valid_1 <= _GEN_195;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1183) begin
                  sectored_entries_5_valid_1 <= _GEN_195;
                end
              end
            end
          end
        end else if (_T_419) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_5_valid_1 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1183) begin
                  sectored_entries_5_valid_1 <= _GEN_195;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1183) begin
                sectored_entries_5_valid_1 <= _GEN_195;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_1 <= _GEN_793;
      end
    end else begin
      sectored_entries_5_valid_1 <= _GEN_523;
    end
    if (_T_3735) begin
      sectored_entries_5_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3104) begin
          if (sectored_entries_5_data_2[0]) begin
            sectored_entries_5_valid_2 <= 1'h0;
          end else if (_T_419) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_5_valid_2 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1183) begin
                    sectored_entries_5_valid_2 <= _GEN_196;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1183) begin
                  sectored_entries_5_valid_2 <= _GEN_196;
                end
              end
            end
          end
        end else if (_T_419) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_5_valid_2 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1183) begin
                  sectored_entries_5_valid_2 <= _GEN_196;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1183) begin
                sectored_entries_5_valid_2 <= _GEN_196;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_2 <= _GEN_794;
      end
    end else begin
      sectored_entries_5_valid_2 <= _GEN_524;
    end
    if (_T_3735) begin
      sectored_entries_5_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3104) begin
          if (sectored_entries_5_data_3[0]) begin
            sectored_entries_5_valid_3 <= 1'h0;
          end else if (_T_419) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_5_valid_3 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1183) begin
                    sectored_entries_5_valid_3 <= _GEN_197;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1183) begin
                  sectored_entries_5_valid_3 <= _GEN_197;
                end
              end
            end
          end
        end else if (_T_419) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_5_valid_3 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1183) begin
                  sectored_entries_5_valid_3 <= _GEN_197;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1183) begin
                sectored_entries_5_valid_3 <= _GEN_197;
              end
            end
          end
        end
      end else begin
        sectored_entries_5_valid_3 <= _GEN_795;
      end
    end else begin
      sectored_entries_5_valid_3 <= _GEN_525;
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1200) begin
            sectored_entries_6_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1200) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_0 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1200) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_1 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1200) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_2 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1200) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_6_data_3 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_3735) begin
      sectored_entries_6_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3251) begin
          if (sectored_entries_6_data_0[0]) begin
            sectored_entries_6_valid_0 <= 1'h0;
          end else if (_T_425) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_6_valid_0 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1200) begin
                    sectored_entries_6_valid_0 <= _GEN_216;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1200) begin
                  sectored_entries_6_valid_0 <= _GEN_216;
                end
              end
            end
          end
        end else if (_T_425) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_6_valid_0 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1200) begin
                  sectored_entries_6_valid_0 <= _GEN_216;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1200) begin
                sectored_entries_6_valid_0 <= _GEN_216;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_0 <= _GEN_820;
      end
    end else begin
      sectored_entries_6_valid_0 <= _GEN_532;
    end
    if (_T_3735) begin
      sectored_entries_6_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3251) begin
          if (sectored_entries_6_data_1[0]) begin
            sectored_entries_6_valid_1 <= 1'h0;
          end else if (_T_425) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_6_valid_1 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1200) begin
                    sectored_entries_6_valid_1 <= _GEN_217;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1200) begin
                  sectored_entries_6_valid_1 <= _GEN_217;
                end
              end
            end
          end
        end else if (_T_425) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_6_valid_1 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1200) begin
                  sectored_entries_6_valid_1 <= _GEN_217;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1200) begin
                sectored_entries_6_valid_1 <= _GEN_217;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_1 <= _GEN_821;
      end
    end else begin
      sectored_entries_6_valid_1 <= _GEN_533;
    end
    if (_T_3735) begin
      sectored_entries_6_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3251) begin
          if (sectored_entries_6_data_2[0]) begin
            sectored_entries_6_valid_2 <= 1'h0;
          end else if (_T_425) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_6_valid_2 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1200) begin
                    sectored_entries_6_valid_2 <= _GEN_218;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1200) begin
                  sectored_entries_6_valid_2 <= _GEN_218;
                end
              end
            end
          end
        end else if (_T_425) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_6_valid_2 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1200) begin
                  sectored_entries_6_valid_2 <= _GEN_218;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1200) begin
                sectored_entries_6_valid_2 <= _GEN_218;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_2 <= _GEN_822;
      end
    end else begin
      sectored_entries_6_valid_2 <= _GEN_534;
    end
    if (_T_3735) begin
      sectored_entries_6_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3251) begin
          if (sectored_entries_6_data_3[0]) begin
            sectored_entries_6_valid_3 <= 1'h0;
          end else if (_T_425) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_6_valid_3 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1200) begin
                    sectored_entries_6_valid_3 <= _GEN_219;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1200) begin
                  sectored_entries_6_valid_3 <= _GEN_219;
                end
              end
            end
          end
        end else if (_T_425) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_6_valid_3 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1200) begin
                  sectored_entries_6_valid_3 <= _GEN_219;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1200) begin
                sectored_entries_6_valid_3 <= _GEN_219;
              end
            end
          end
        end
      end else begin
        sectored_entries_6_valid_3 <= _GEN_823;
      end
    end else begin
      sectored_entries_6_valid_3 <= _GEN_535;
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1217) begin
            sectored_entries_7_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1217) begin
            if (2'h0 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_0 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1217) begin
            if (2'h1 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_1 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1217) begin
            if (2'h2 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_2 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (!(_T_1032)) begin
          if (_T_1217) begin
            if (2'h3 == r_refill_tag[1:0]) begin
              sectored_entries_7_data_3 <= _T_1031;
            end
          end
        end
      end
    end
    if (_T_3735) begin
      sectored_entries_7_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3398) begin
          if (sectored_entries_7_data_0[0]) begin
            sectored_entries_7_valid_0 <= 1'h0;
          end else if (_T_431) begin
            if (2'h0 == vpn[1:0]) begin
              sectored_entries_7_valid_0 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1217) begin
                    sectored_entries_7_valid_0 <= _GEN_238;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1217) begin
                  sectored_entries_7_valid_0 <= _GEN_238;
                end
              end
            end
          end
        end else if (_T_431) begin
          if (2'h0 == vpn[1:0]) begin
            sectored_entries_7_valid_0 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1217) begin
                  sectored_entries_7_valid_0 <= _GEN_238;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1217) begin
                sectored_entries_7_valid_0 <= _GEN_238;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_0 <= _GEN_848;
      end
    end else begin
      sectored_entries_7_valid_0 <= _GEN_542;
    end
    if (_T_3735) begin
      sectored_entries_7_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3398) begin
          if (sectored_entries_7_data_1[0]) begin
            sectored_entries_7_valid_1 <= 1'h0;
          end else if (_T_431) begin
            if (2'h1 == vpn[1:0]) begin
              sectored_entries_7_valid_1 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1217) begin
                    sectored_entries_7_valid_1 <= _GEN_239;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1217) begin
                  sectored_entries_7_valid_1 <= _GEN_239;
                end
              end
            end
          end
        end else if (_T_431) begin
          if (2'h1 == vpn[1:0]) begin
            sectored_entries_7_valid_1 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1217) begin
                  sectored_entries_7_valid_1 <= _GEN_239;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1217) begin
                sectored_entries_7_valid_1 <= _GEN_239;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_1 <= _GEN_849;
      end
    end else begin
      sectored_entries_7_valid_1 <= _GEN_543;
    end
    if (_T_3735) begin
      sectored_entries_7_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3398) begin
          if (sectored_entries_7_data_2[0]) begin
            sectored_entries_7_valid_2 <= 1'h0;
          end else if (_T_431) begin
            if (2'h2 == vpn[1:0]) begin
              sectored_entries_7_valid_2 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1217) begin
                    sectored_entries_7_valid_2 <= _GEN_240;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1217) begin
                  sectored_entries_7_valid_2 <= _GEN_240;
                end
              end
            end
          end
        end else if (_T_431) begin
          if (2'h2 == vpn[1:0]) begin
            sectored_entries_7_valid_2 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1217) begin
                  sectored_entries_7_valid_2 <= _GEN_240;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1217) begin
                sectored_entries_7_valid_2 <= _GEN_240;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_2 <= _GEN_850;
      end
    end else begin
      sectored_entries_7_valid_2 <= _GEN_544;
    end
    if (_T_3735) begin
      sectored_entries_7_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_3398) begin
          if (sectored_entries_7_data_3[0]) begin
            sectored_entries_7_valid_3 <= 1'h0;
          end else if (_T_431) begin
            if (2'h3 == vpn[1:0]) begin
              sectored_entries_7_valid_3 <= 1'h0;
            end else if (_T_993) begin
              if (!(_T_1015)) begin
                if (!(_T_1032)) begin
                  if (_T_1217) begin
                    sectored_entries_7_valid_3 <= _GEN_241;
                  end
                end
              end
            end
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1217) begin
                  sectored_entries_7_valid_3 <= _GEN_241;
                end
              end
            end
          end
        end else if (_T_431) begin
          if (2'h3 == vpn[1:0]) begin
            sectored_entries_7_valid_3 <= 1'h0;
          end else if (_T_993) begin
            if (!(_T_1015)) begin
              if (!(_T_1032)) begin
                if (_T_1217) begin
                  sectored_entries_7_valid_3 <= _GEN_241;
                end
              end
            end
          end
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (!(_T_1032)) begin
              if (_T_1217) begin
                sectored_entries_7_valid_3 <= _GEN_241;
              end
            end
          end
        end
      end else begin
        sectored_entries_7_valid_3 <= _GEN_851;
      end
    end else begin
      sectored_entries_7_valid_3 <= _GEN_545;
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          if (_T_1033) begin
            superpage_entries_0_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          if (_T_1033) begin
            superpage_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          if (_T_1033) begin
            superpage_entries_0_data_0 <= _T_1031;
          end
        end
      end
    end
    if (_T_3735) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_0) begin
          superpage_entries_0_valid_0 <= 1'h0;
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (_T_1032) begin
              superpage_entries_0_valid_0 <= _GEN_66;
            end
          end
        end
      end else begin
        superpage_entries_0_valid_0 <= _GEN_858;
      end
    end else if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          superpage_entries_0_valid_0 <= _GEN_66;
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          if (_T_1049) begin
            superpage_entries_1_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          if (_T_1049) begin
            superpage_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          if (_T_1049) begin
            superpage_entries_1_data_0 <= _T_1031;
          end
        end
      end
    end
    if (_T_3735) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_1) begin
          superpage_entries_1_valid_0 <= 1'h0;
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (_T_1032) begin
              superpage_entries_1_valid_0 <= _GEN_70;
            end
          end
        end
      end else begin
        superpage_entries_1_valid_0 <= _GEN_862;
      end
    end else if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          superpage_entries_1_valid_0 <= _GEN_70;
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          if (_T_1065) begin
            superpage_entries_2_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          if (_T_1065) begin
            superpage_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          if (_T_1065) begin
            superpage_entries_2_data_0 <= _T_1031;
          end
        end
      end
    end
    if (_T_3735) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_2) begin
          superpage_entries_2_valid_0 <= 1'h0;
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (_T_1032) begin
              superpage_entries_2_valid_0 <= _GEN_74;
            end
          end
        end
      end else begin
        superpage_entries_2_valid_0 <= _GEN_866;
      end
    end else if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          superpage_entries_2_valid_0 <= _GEN_74;
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          if (_T_1081) begin
            superpage_entries_3_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          if (_T_1081) begin
            superpage_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          if (_T_1081) begin
            superpage_entries_3_data_0 <= _T_1031;
          end
        end
      end
    end
    if (_T_3735) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_3) begin
          superpage_entries_3_valid_0 <= 1'h0;
        end else if (_T_993) begin
          if (!(_T_1015)) begin
            if (_T_1032) begin
              superpage_entries_3_valid_0 <= _GEN_78;
            end
          end
        end
      end else begin
        superpage_entries_3_valid_0 <= _GEN_870;
      end
    end else if (_T_993) begin
      if (!(_T_1015)) begin
        if (_T_1032) begin
          superpage_entries_3_valid_0 <= _GEN_78;
        end
      end
    end
    if (_T_993) begin
      if (_T_1015) begin
        special_entry_level <= io_ptw_resp_bits_level;
      end
    end
    if (_T_993) begin
      if (_T_1015) begin
        special_entry_tag <= r_refill_tag;
      end
    end
    if (_T_993) begin
      if (_T_1015) begin
        special_entry_data_0 <= _T_1031;
      end
    end
    if (_T_3735) begin
      special_entry_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_656) begin
          special_entry_valid_0 <= 1'h0;
        end else if (_T_993) begin
          special_entry_valid_0 <= _GEN_354;
        end
      end else begin
        special_entry_valid_0 <= _GEN_874;
      end
    end else if (_T_993) begin
      special_entry_valid_0 <= _GEN_354;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if (_T_2355) begin
      state <= 2'h3;
    end else if (_T_4) begin
      if (io_kill) begin
        state <= 2'h0;
      end else if (io_ptw_req_ready) begin
        if (io_sfence_valid) begin
          state <= 2'h3;
        end else begin
          state <= 2'h2;
        end
      end else if (io_sfence_valid) begin
        state <= 2'h0;
      end else if (_T_2225) begin
        state <= 2'h1;
      end
    end else if (_T_2225) begin
      state <= 2'h1;
    end
    if (_T_2225) begin
      r_refill_tag <= vpn;
    end
    if (_T_2225) begin
      if (_T_2245) begin
        r_superpage_repl_addr <= _T_2240[1:0];
      end else if (_T_2246[0]) begin
        r_superpage_repl_addr <= 2'h0;
      end else if (_T_2246[1]) begin
        r_superpage_repl_addr <= 2'h1;
      end else if (_T_2246[2]) begin
        r_superpage_repl_addr <= 2'h2;
      end else begin
        r_superpage_repl_addr <= 2'h3;
      end
    end
    if (_T_2225) begin
      if (_T_2309) begin
        r_sectored_repl_addr <= _T_2276[2:0];
      end else if (_T_2310[0]) begin
        r_sectored_repl_addr <= 3'h0;
      end else if (_T_2310[1]) begin
        r_sectored_repl_addr <= 3'h1;
      end else if (_T_2310[2]) begin
        r_sectored_repl_addr <= 3'h2;
      end else if (_T_2310[3]) begin
        r_sectored_repl_addr <= 3'h3;
      end else if (_T_2310[4]) begin
        r_sectored_repl_addr <= 3'h4;
      end else if (_T_2310[5]) begin
        r_sectored_repl_addr <= 3'h5;
      end else if (_T_2310[6]) begin
        r_sectored_repl_addr <= 3'h6;
      end else begin
        r_sectored_repl_addr <= 3'h7;
      end
    end
    if (_T_2225) begin
      r_sectored_hit_addr <= _T_2042;
    end
    if (_T_2225) begin
      r_sectored_hit <= _T_2024;
    end
    if (_T_2017) begin
      if (_T_2024) begin
        _T_2015 <= _T_2069[7:1];
      end
    end
    if (_T_2017) begin
      if (_T_2074) begin
        _T_2016 <= _T_2101[3:1];
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & _T_2362) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:368 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"); // @[TLB.scala 368:13:chipyard.TestHarness.RocketConfig.fir@224425.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_sfence_valid & _T_2362) begin
          $fatal; // @[TLB.scala 368:13:chipyard.TestHarness.RocketConfig.fir@224426.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
