module TLMonitor_41( // @[:chipyard.TestHarness.RocketConfig.fir@102456.2]
  input         clock, // @[:chipyard.TestHarness.RocketConfig.fir@102457.4]
  input         reset, // @[:chipyard.TestHarness.RocketConfig.fir@102458.4]
  input         io_in_a_ready, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input         io_in_a_valid, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [2:0]  io_in_a_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [2:0]  io_in_a_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [2:0]  io_in_a_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [2:0]  io_in_a_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [31:0] io_in_a_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [7:0]  io_in_a_bits_mask, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input         io_in_a_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input         io_in_b_ready, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input         io_in_b_valid, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [1:0]  io_in_b_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [31:0] io_in_b_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input         io_in_c_ready, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input         io_in_c_valid, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [2:0]  io_in_c_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [2:0]  io_in_c_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [2:0]  io_in_c_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [2:0]  io_in_c_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [31:0] io_in_c_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input         io_in_c_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input         io_in_d_ready, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input         io_in_d_valid, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [2:0]  io_in_d_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [1:0]  io_in_d_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [2:0]  io_in_d_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [2:0]  io_in_d_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [2:0]  io_in_d_bits_sink, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input         io_in_d_bits_denied, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input         io_in_d_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input         io_in_e_valid, // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
  input  [2:0]  io_in_e_bits_sink // @[:chipyard.TestHarness.RocketConfig.fir@102459.4]
);
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104949.4]
  wire  _T_4; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@102470.6]
  wire  _T_5; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@102471.6]
  wire  _T_6; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@102472.6]
  wire  _T_7; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@102473.6]
  wire  _T_9; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@102480.6]
  wire  _T_10; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@102481.6]
  wire  _T_11; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@102482.6]
  wire [12:0] _T_13; // @[package.scala 189:77:chipyard.TestHarness.RocketConfig.fir@102484.6]
  wire [5:0] _T_15; // @[package.scala 189:46:chipyard.TestHarness.RocketConfig.fir@102486.6]
  wire [31:0] _GEN_71; // @[Edges.scala 22:16:chipyard.TestHarness.RocketConfig.fir@102487.6]
  wire [31:0] _T_16; // @[Edges.scala 22:16:chipyard.TestHarness.RocketConfig.fir@102487.6]
  wire  _T_17; // @[Edges.scala 22:24:chipyard.TestHarness.RocketConfig.fir@102488.6]
  wire [3:0] _T_20; // @[OneHot.scala 65:12:chipyard.TestHarness.RocketConfig.fir@102491.6]
  wire [2:0] _T_22; // @[Misc.scala 201:81:chipyard.TestHarness.RocketConfig.fir@102493.6]
  wire  _T_23; // @[Misc.scala 205:21:chipyard.TestHarness.RocketConfig.fir@102494.6]
  wire  _T_26; // @[Misc.scala 210:20:chipyard.TestHarness.RocketConfig.fir@102497.6]
  wire  _T_28; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102499.6]
  wire  _T_29; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102500.6]
  wire  _T_31; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102502.6]
  wire  _T_32; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102503.6]
  wire  _T_35; // @[Misc.scala 210:20:chipyard.TestHarness.RocketConfig.fir@102506.6]
  wire  _T_36; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102507.6]
  wire  _T_37; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102508.6]
  wire  _T_38; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102509.6]
  wire  _T_39; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102510.6]
  wire  _T_40; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102511.6]
  wire  _T_41; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102512.6]
  wire  _T_42; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102513.6]
  wire  _T_43; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102514.6]
  wire  _T_44; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102515.6]
  wire  _T_45; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102516.6]
  wire  _T_46; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102517.6]
  wire  _T_47; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102518.6]
  wire  _T_50; // @[Misc.scala 210:20:chipyard.TestHarness.RocketConfig.fir@102521.6]
  wire  _T_51; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102522.6]
  wire  _T_52; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102523.6]
  wire  _T_53; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102524.6]
  wire  _T_54; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102525.6]
  wire  _T_55; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102526.6]
  wire  _T_56; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102527.6]
  wire  _T_57; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102528.6]
  wire  _T_58; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102529.6]
  wire  _T_59; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102530.6]
  wire  _T_60; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102531.6]
  wire  _T_61; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102532.6]
  wire  _T_62; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102533.6]
  wire  _T_63; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102534.6]
  wire  _T_64; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102535.6]
  wire  _T_65; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102536.6]
  wire  _T_66; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102537.6]
  wire  _T_67; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102538.6]
  wire  _T_68; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102539.6]
  wire  _T_69; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102540.6]
  wire  _T_70; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102541.6]
  wire  _T_71; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102542.6]
  wire  _T_72; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102543.6]
  wire  _T_73; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102544.6]
  wire  _T_74; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102545.6]
  wire [7:0] _T_81; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@102552.6]
  wire  _T_120; // @[Monitor.scala 79:25:chipyard.TestHarness.RocketConfig.fir@102595.6]
  wire  _T_121; // @[Parameters.scala 92:48:chipyard.TestHarness.RocketConfig.fir@102597.8]
  wire [31:0] _T_123; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@102599.8]
  wire [32:0] _T_124; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@102600.8]
  wire [32:0] _T_126; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@102602.8]
  wire  _T_127; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@102603.8]
  wire  _T_128; // @[Parameters.scala 551:56:chipyard.TestHarness.RocketConfig.fir@102604.8]
  wire  _T_131; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102607.8]
  wire  _T_132; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102608.8]
  wire  _T_140; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@102625.8]
  wire  _T_148; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102634.8]
  wire  _T_149; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102635.8]
  wire  _T_151; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102641.8]
  wire  _T_152; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102642.8]
  wire  _T_155; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102649.8]
  wire  _T_156; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102650.8]
  wire  _T_158; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102656.8]
  wire  _T_159; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102657.8]
  wire  _T_160; // @[Bundles.scala 110:27:chipyard.TestHarness.RocketConfig.fir@102662.8]
  wire  _T_162; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102664.8]
  wire  _T_163; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102665.8]
  wire [7:0] _T_164; // @[Monitor.scala 86:18:chipyard.TestHarness.RocketConfig.fir@102670.8]
  wire  _T_165; // @[Monitor.scala 86:31:chipyard.TestHarness.RocketConfig.fir@102671.8]
  wire  _T_167; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102673.8]
  wire  _T_168; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102674.8]
  wire  _T_169; // @[Monitor.scala 87:18:chipyard.TestHarness.RocketConfig.fir@102679.8]
  wire  _T_171; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102681.8]
  wire  _T_172; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102682.8]
  wire  _T_173; // @[Monitor.scala 90:25:chipyard.TestHarness.RocketConfig.fir@102688.6]
  wire  _T_217; // @[Monitor.scala 97:31:chipyard.TestHarness.RocketConfig.fir@102763.8]
  wire  _T_219; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102765.8]
  wire  _T_220; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102766.8]
  wire  _T_230; // @[Monitor.scala 102:25:chipyard.TestHarness.RocketConfig.fir@102789.6]
  wire  _T_232; // @[Parameters.scala 93:42:chipyard.TestHarness.RocketConfig.fir@102792.8]
  wire  _T_240; // @[Parameters.scala 551:56:chipyard.TestHarness.RocketConfig.fir@102800.8]
  wire  _T_243; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102803.8]
  wire  _T_244; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102804.8]
  wire  _T_251; // @[Monitor.scala 106:31:chipyard.TestHarness.RocketConfig.fir@102823.8]
  wire  _T_253; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102825.8]
  wire  _T_254; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102826.8]
  wire  _T_255; // @[Monitor.scala 107:30:chipyard.TestHarness.RocketConfig.fir@102831.8]
  wire  _T_257; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102833.8]
  wire  _T_258; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102834.8]
  wire  _T_263; // @[Monitor.scala 111:25:chipyard.TestHarness.RocketConfig.fir@102848.6]
  wire  _T_292; // @[Monitor.scala 119:25:chipyard.TestHarness.RocketConfig.fir@102899.6]
  wire [7:0] _T_317; // @[Monitor.scala 124:33:chipyard.TestHarness.RocketConfig.fir@102941.8]
  wire [7:0] _T_318; // @[Monitor.scala 124:31:chipyard.TestHarness.RocketConfig.fir@102942.8]
  wire  _T_319; // @[Monitor.scala 124:40:chipyard.TestHarness.RocketConfig.fir@102943.8]
  wire  _T_321; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102945.8]
  wire  _T_322; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102946.8]
  wire  _T_323; // @[Monitor.scala 127:25:chipyard.TestHarness.RocketConfig.fir@102952.6]
  wire  _T_325; // @[Parameters.scala 93:42:chipyard.TestHarness.RocketConfig.fir@102955.8]
  wire  _T_333; // @[Parameters.scala 551:56:chipyard.TestHarness.RocketConfig.fir@102963.8]
  wire  _T_336; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102966.8]
  wire  _T_337; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102967.8]
  wire  _T_344; // @[Bundles.scala 140:33:chipyard.TestHarness.RocketConfig.fir@102986.8]
  wire  _T_346; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102988.8]
  wire  _T_347; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102989.8]
  wire  _T_352; // @[Monitor.scala 135:25:chipyard.TestHarness.RocketConfig.fir@103003.6]
  wire  _T_373; // @[Bundles.scala 147:30:chipyard.TestHarness.RocketConfig.fir@103037.8]
  wire  _T_375; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103039.8]
  wire  _T_376; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103040.8]
  wire  _T_381; // @[Monitor.scala 143:25:chipyard.TestHarness.RocketConfig.fir@103054.6]
  wire  _T_402; // @[Bundles.scala 160:28:chipyard.TestHarness.RocketConfig.fir@103088.8]
  wire  _T_404; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103090.8]
  wire  _T_405; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103091.8]
  wire  _T_414; // @[Bundles.scala 44:24:chipyard.TestHarness.RocketConfig.fir@103115.6]
  wire  _T_416; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103117.6]
  wire  _T_417; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103118.6]
  wire  _T_418; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103123.6]
  wire  _T_419; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103124.6]
  wire  _T_420; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103125.6]
  wire  _T_421; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103126.6]
  wire  _T_423; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@103133.6]
  wire  _T_424; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@103134.6]
  wire  _T_425; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@103135.6]
  wire  _T_426; // @[Monitor.scala 303:31:chipyard.TestHarness.RocketConfig.fir@103136.6]
  wire  _T_427; // @[Monitor.scala 307:25:chipyard.TestHarness.RocketConfig.fir@103137.6]
  wire  _T_429; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103140.8]
  wire  _T_430; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103141.8]
  wire  _T_431; // @[Monitor.scala 309:27:chipyard.TestHarness.RocketConfig.fir@103146.8]
  wire  _T_433; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103148.8]
  wire  _T_434; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103149.8]
  wire  _T_435; // @[Monitor.scala 310:28:chipyard.TestHarness.RocketConfig.fir@103154.8]
  wire  _T_437; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103156.8]
  wire  _T_438; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103157.8]
  wire  _T_439; // @[Monitor.scala 311:15:chipyard.TestHarness.RocketConfig.fir@103162.8]
  wire  _T_441; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103164.8]
  wire  _T_442; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103165.8]
  wire  _T_443; // @[Monitor.scala 312:15:chipyard.TestHarness.RocketConfig.fir@103170.8]
  wire  _T_445; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103172.8]
  wire  _T_446; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103173.8]
  wire  _T_447; // @[Monitor.scala 315:25:chipyard.TestHarness.RocketConfig.fir@103179.6]
  wire  _T_452; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103189.8]
  wire  _T_453; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103190.8]
  wire  _T_458; // @[Bundles.scala 104:26:chipyard.TestHarness.RocketConfig.fir@103203.8]
  wire  _T_460; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103205.8]
  wire  _T_461; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103206.8]
  wire  _T_462; // @[Monitor.scala 320:28:chipyard.TestHarness.RocketConfig.fir@103211.8]
  wire  _T_464; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103213.8]
  wire  _T_465; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103214.8]
  wire  _T_475; // @[Monitor.scala 325:25:chipyard.TestHarness.RocketConfig.fir@103237.6]
  wire  _T_495; // @[Monitor.scala 331:30:chipyard.TestHarness.RocketConfig.fir@103278.8]
  wire  _T_497; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103280.8]
  wire  _T_498; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103281.8]
  wire  _T_504; // @[Monitor.scala 335:25:chipyard.TestHarness.RocketConfig.fir@103296.6]
  wire  _T_521; // @[Monitor.scala 343:25:chipyard.TestHarness.RocketConfig.fir@103331.6]
  wire  _T_539; // @[Monitor.scala 351:25:chipyard.TestHarness.RocketConfig.fir@103367.6]
  wire [31:0] _T_598; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@103454.6]
  wire [32:0] _T_599; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@103455.6]
  wire [32:0] _T_601; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@103457.6]
  wire  _T_602; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@103458.6]
  wire [31:0] _T_608; // @[Edges.scala 22:16:chipyard.TestHarness.RocketConfig.fir@103466.6]
  wire  _T_609; // @[Edges.scala 22:24:chipyard.TestHarness.RocketConfig.fir@103467.6]
  wire  _T_707; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103582.8]
  wire  _T_708; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103583.8]
  wire  _T_713; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103596.8]
  wire  _T_714; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103597.8]
  wire  _T_715; // @[Bundles.scala 104:26:chipyard.TestHarness.RocketConfig.fir@103602.8]
  wire  _T_717; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103604.8]
  wire  _T_718; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103605.8]
  wire  _T_863; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103929.6]
  wire  _T_864; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103930.6]
  wire  _T_865; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103931.6]
  wire  _T_866; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103932.6]
  wire  _T_868; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@103939.6]
  wire  _T_869; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@103940.6]
  wire  _T_870; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@103941.6]
  wire [12:0] _T_872; // @[package.scala 189:77:chipyard.TestHarness.RocketConfig.fir@103943.6]
  wire [5:0] _T_874; // @[package.scala 189:46:chipyard.TestHarness.RocketConfig.fir@103945.6]
  wire [31:0] _GEN_72; // @[Edges.scala 22:16:chipyard.TestHarness.RocketConfig.fir@103946.6]
  wire [31:0] _T_875; // @[Edges.scala 22:16:chipyard.TestHarness.RocketConfig.fir@103946.6]
  wire  _T_876; // @[Edges.scala 22:24:chipyard.TestHarness.RocketConfig.fir@103947.6]
  wire [31:0] _T_877; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@103948.6]
  wire [32:0] _T_878; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@103949.6]
  wire [32:0] _T_880; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@103951.6]
  wire  _T_881; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@103952.6]
  wire  _T_921; // @[Monitor.scala 239:25:chipyard.TestHarness.RocketConfig.fir@103998.6]
  wire  _T_923; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104001.8]
  wire  _T_924; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104002.8]
  wire  _T_926; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104008.8]
  wire  _T_927; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104009.8]
  wire  _T_928; // @[Monitor.scala 242:30:chipyard.TestHarness.RocketConfig.fir@104014.8]
  wire  _T_930; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104016.8]
  wire  _T_931; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104017.8]
  wire  _T_933; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104023.8]
  wire  _T_934; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104024.8]
  wire  _T_935; // @[Bundles.scala 122:29:chipyard.TestHarness.RocketConfig.fir@104029.8]
  wire  _T_937; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104031.8]
  wire  _T_938; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104032.8]
  wire  _T_939; // @[Monitor.scala 245:18:chipyard.TestHarness.RocketConfig.fir@104037.8]
  wire  _T_941; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104039.8]
  wire  _T_942; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104040.8]
  wire  _T_943; // @[Monitor.scala 248:25:chipyard.TestHarness.RocketConfig.fir@104046.6]
  wire  _T_961; // @[Monitor.scala 256:25:chipyard.TestHarness.RocketConfig.fir@104086.6]
  wire  _T_962; // @[Parameters.scala 92:48:chipyard.TestHarness.RocketConfig.fir@104088.8]
  wire  _T_969; // @[Parameters.scala 551:56:chipyard.TestHarness.RocketConfig.fir@104095.8]
  wire  _T_972; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104098.8]
  wire  _T_973; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104099.8]
  wire  _T_981; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@104116.8]
  wire  _T_989; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104125.8]
  wire  _T_990; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104126.8]
  wire  _T_1001; // @[Bundles.scala 116:29:chipyard.TestHarness.RocketConfig.fir@104153.8]
  wire  _T_1003; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104155.8]
  wire  _T_1004; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104156.8]
  wire  _T_1009; // @[Monitor.scala 266:25:chipyard.TestHarness.RocketConfig.fir@104170.6]
  wire  _T_1053; // @[Monitor.scala 275:25:chipyard.TestHarness.RocketConfig.fir@104246.6]
  wire  _T_1063; // @[Monitor.scala 279:31:chipyard.TestHarness.RocketConfig.fir@104269.8]
  wire  _T_1065; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104271.8]
  wire  _T_1066; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104272.8]
  wire  _T_1071; // @[Monitor.scala 283:25:chipyard.TestHarness.RocketConfig.fir@104286.6]
  wire  _T_1085; // @[Monitor.scala 290:25:chipyard.TestHarness.RocketConfig.fir@104318.6]
  wire  _T_1103; // @[Monitor.scala 361:31:chipyard.TestHarness.RocketConfig.fir@104360.6]
  wire  _T_1105; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104362.6]
  wire  _T_1106; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104363.6]
  wire  _T_1107; // @[Decoupled.scala 40:37:chipyard.TestHarness.RocketConfig.fir@104369.4]
  wire  _T_1114; // @[Edges.scala 93:28:chipyard.TestHarness.RocketConfig.fir@104376.4]
  reg [2:0] _T_1116; // @[Edges.scala 230:27:chipyard.TestHarness.RocketConfig.fir@104378.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_1118; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104380.4]
  wire  _T_1119; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104381.4]
  reg [2:0] _T_1127; // @[Monitor.scala 381:22:chipyard.TestHarness.RocketConfig.fir@104392.4]
  reg [31:0] _RAND_1;
  reg [2:0] _T_1128; // @[Monitor.scala 382:22:chipyard.TestHarness.RocketConfig.fir@104393.4]
  reg [31:0] _RAND_2;
  reg [2:0] _T_1129; // @[Monitor.scala 383:22:chipyard.TestHarness.RocketConfig.fir@104394.4]
  reg [31:0] _RAND_3;
  reg [2:0] _T_1130; // @[Monitor.scala 384:22:chipyard.TestHarness.RocketConfig.fir@104395.4]
  reg [31:0] _RAND_4;
  reg [31:0] _T_1131; // @[Monitor.scala 385:22:chipyard.TestHarness.RocketConfig.fir@104396.4]
  reg [31:0] _RAND_5;
  wire  _T_1132; // @[Monitor.scala 386:22:chipyard.TestHarness.RocketConfig.fir@104397.4]
  wire  _T_1133; // @[Monitor.scala 386:19:chipyard.TestHarness.RocketConfig.fir@104398.4]
  wire  _T_1134; // @[Monitor.scala 387:32:chipyard.TestHarness.RocketConfig.fir@104400.6]
  wire  _T_1136; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104402.6]
  wire  _T_1137; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104403.6]
  wire  _T_1138; // @[Monitor.scala 388:32:chipyard.TestHarness.RocketConfig.fir@104408.6]
  wire  _T_1140; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104410.6]
  wire  _T_1141; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104411.6]
  wire  _T_1142; // @[Monitor.scala 389:32:chipyard.TestHarness.RocketConfig.fir@104416.6]
  wire  _T_1144; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104418.6]
  wire  _T_1145; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104419.6]
  wire  _T_1146; // @[Monitor.scala 390:32:chipyard.TestHarness.RocketConfig.fir@104424.6]
  wire  _T_1148; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104426.6]
  wire  _T_1149; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104427.6]
  wire  _T_1150; // @[Monitor.scala 391:32:chipyard.TestHarness.RocketConfig.fir@104432.6]
  wire  _T_1152; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104434.6]
  wire  _T_1153; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104435.6]
  wire  _T_1155; // @[Monitor.scala 393:20:chipyard.TestHarness.RocketConfig.fir@104442.4]
  wire  _T_1156; // @[Decoupled.scala 40:37:chipyard.TestHarness.RocketConfig.fir@104450.4]
  wire [12:0] _T_1158; // @[package.scala 189:77:chipyard.TestHarness.RocketConfig.fir@104452.4]
  wire [5:0] _T_1160; // @[package.scala 189:46:chipyard.TestHarness.RocketConfig.fir@104454.4]
  reg [2:0] _T_1164; // @[Edges.scala 230:27:chipyard.TestHarness.RocketConfig.fir@104458.4]
  reg [31:0] _RAND_6;
  wire [2:0] _T_1166; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104460.4]
  wire  _T_1167; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104461.4]
  reg [2:0] _T_1175; // @[Monitor.scala 532:22:chipyard.TestHarness.RocketConfig.fir@104472.4]
  reg [31:0] _RAND_7;
  reg [1:0] _T_1176; // @[Monitor.scala 533:22:chipyard.TestHarness.RocketConfig.fir@104473.4]
  reg [31:0] _RAND_8;
  reg [2:0] _T_1177; // @[Monitor.scala 534:22:chipyard.TestHarness.RocketConfig.fir@104474.4]
  reg [31:0] _RAND_9;
  reg [2:0] _T_1178; // @[Monitor.scala 535:22:chipyard.TestHarness.RocketConfig.fir@104475.4]
  reg [31:0] _RAND_10;
  reg [2:0] _T_1179; // @[Monitor.scala 536:22:chipyard.TestHarness.RocketConfig.fir@104476.4]
  reg [31:0] _RAND_11;
  reg  _T_1180; // @[Monitor.scala 537:22:chipyard.TestHarness.RocketConfig.fir@104477.4]
  reg [31:0] _RAND_12;
  wire  _T_1181; // @[Monitor.scala 538:22:chipyard.TestHarness.RocketConfig.fir@104478.4]
  wire  _T_1182; // @[Monitor.scala 538:19:chipyard.TestHarness.RocketConfig.fir@104479.4]
  wire  _T_1183; // @[Monitor.scala 539:29:chipyard.TestHarness.RocketConfig.fir@104481.6]
  wire  _T_1185; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104483.6]
  wire  _T_1186; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104484.6]
  wire  _T_1187; // @[Monitor.scala 540:29:chipyard.TestHarness.RocketConfig.fir@104489.6]
  wire  _T_1189; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104491.6]
  wire  _T_1190; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104492.6]
  wire  _T_1191; // @[Monitor.scala 541:29:chipyard.TestHarness.RocketConfig.fir@104497.6]
  wire  _T_1193; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104499.6]
  wire  _T_1194; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104500.6]
  wire  _T_1195; // @[Monitor.scala 542:29:chipyard.TestHarness.RocketConfig.fir@104505.6]
  wire  _T_1197; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104507.6]
  wire  _T_1198; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104508.6]
  wire  _T_1199; // @[Monitor.scala 543:29:chipyard.TestHarness.RocketConfig.fir@104513.6]
  wire  _T_1201; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104515.6]
  wire  _T_1202; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104516.6]
  wire  _T_1203; // @[Monitor.scala 544:29:chipyard.TestHarness.RocketConfig.fir@104521.6]
  wire  _T_1205; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104523.6]
  wire  _T_1206; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104524.6]
  wire  _T_1208; // @[Monitor.scala 546:20:chipyard.TestHarness.RocketConfig.fir@104531.4]
  wire  _T_1209; // @[Decoupled.scala 40:37:chipyard.TestHarness.RocketConfig.fir@104540.4]
  reg [2:0] _T_1218; // @[Edges.scala 230:27:chipyard.TestHarness.RocketConfig.fir@104549.4]
  reg [31:0] _RAND_13;
  wire [2:0] _T_1220; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104551.4]
  wire  _T_1221; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104552.4]
  reg [1:0] _T_1230; // @[Monitor.scala 405:22:chipyard.TestHarness.RocketConfig.fir@104564.4]
  reg [31:0] _RAND_14;
  reg [31:0] _T_1233; // @[Monitor.scala 408:22:chipyard.TestHarness.RocketConfig.fir@104567.4]
  reg [31:0] _RAND_15;
  wire  _T_1234; // @[Monitor.scala 409:22:chipyard.TestHarness.RocketConfig.fir@104568.4]
  wire  _T_1235; // @[Monitor.scala 409:19:chipyard.TestHarness.RocketConfig.fir@104569.4]
  wire  _T_1240; // @[Monitor.scala 411:32:chipyard.TestHarness.RocketConfig.fir@104579.6]
  wire  _T_1242; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104581.6]
  wire  _T_1243; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104582.6]
  wire  _T_1252; // @[Monitor.scala 414:32:chipyard.TestHarness.RocketConfig.fir@104603.6]
  wire  _T_1254; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104605.6]
  wire  _T_1255; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104606.6]
  wire  _T_1257; // @[Monitor.scala 416:20:chipyard.TestHarness.RocketConfig.fir@104613.4]
  wire  _T_1258; // @[Decoupled.scala 40:37:chipyard.TestHarness.RocketConfig.fir@104621.4]
  reg [2:0] _T_1266; // @[Edges.scala 230:27:chipyard.TestHarness.RocketConfig.fir@104629.4]
  reg [31:0] _RAND_16;
  wire [2:0] _T_1268; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104631.4]
  wire  _T_1269; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104632.4]
  reg [2:0] _T_1277; // @[Monitor.scala 509:22:chipyard.TestHarness.RocketConfig.fir@104643.4]
  reg [31:0] _RAND_17;
  reg [2:0] _T_1278; // @[Monitor.scala 510:22:chipyard.TestHarness.RocketConfig.fir@104644.4]
  reg [31:0] _RAND_18;
  reg [2:0] _T_1279; // @[Monitor.scala 511:22:chipyard.TestHarness.RocketConfig.fir@104645.4]
  reg [31:0] _RAND_19;
  reg [2:0] _T_1280; // @[Monitor.scala 512:22:chipyard.TestHarness.RocketConfig.fir@104646.4]
  reg [31:0] _RAND_20;
  reg [31:0] _T_1281; // @[Monitor.scala 513:22:chipyard.TestHarness.RocketConfig.fir@104647.4]
  reg [31:0] _RAND_21;
  wire  _T_1282; // @[Monitor.scala 514:22:chipyard.TestHarness.RocketConfig.fir@104648.4]
  wire  _T_1283; // @[Monitor.scala 514:19:chipyard.TestHarness.RocketConfig.fir@104649.4]
  wire  _T_1284; // @[Monitor.scala 515:32:chipyard.TestHarness.RocketConfig.fir@104651.6]
  wire  _T_1286; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104653.6]
  wire  _T_1287; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104654.6]
  wire  _T_1288; // @[Monitor.scala 516:32:chipyard.TestHarness.RocketConfig.fir@104659.6]
  wire  _T_1290; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104661.6]
  wire  _T_1291; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104662.6]
  wire  _T_1292; // @[Monitor.scala 517:32:chipyard.TestHarness.RocketConfig.fir@104667.6]
  wire  _T_1294; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104669.6]
  wire  _T_1295; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104670.6]
  wire  _T_1296; // @[Monitor.scala 518:32:chipyard.TestHarness.RocketConfig.fir@104675.6]
  wire  _T_1298; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104677.6]
  wire  _T_1299; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104678.6]
  wire  _T_1300; // @[Monitor.scala 519:32:chipyard.TestHarness.RocketConfig.fir@104683.6]
  wire  _T_1302; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104685.6]
  wire  _T_1303; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104686.6]
  wire  _T_1305; // @[Monitor.scala 521:20:chipyard.TestHarness.RocketConfig.fir@104693.4]
  reg [4:0] inflight; // @[Monitor.scala 608:27:chipyard.TestHarness.RocketConfig.fir@104701.4]
  reg [31:0] _RAND_22;
  reg [19:0] inflight_opcodes; // @[Monitor.scala 610:35:chipyard.TestHarness.RocketConfig.fir@104702.4]
  reg [31:0] _RAND_23;
  reg [19:0] inflight_sizes; // @[Monitor.scala 612:33:chipyard.TestHarness.RocketConfig.fir@104703.4]
  reg [31:0] _RAND_24;
  reg [2:0] _T_1315; // @[Edges.scala 230:27:chipyard.TestHarness.RocketConfig.fir@104713.4]
  reg [31:0] _RAND_25;
  wire [2:0] _T_1317; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104715.4]
  wire  a_first; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104716.4]
  reg [2:0] _T_1333; // @[Edges.scala 230:27:chipyard.TestHarness.RocketConfig.fir@104735.4]
  reg [31:0] _RAND_26;
  wire [2:0] _T_1335; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104737.4]
  wire  d_first; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104738.4]
  wire [4:0] _GEN_73; // @[Monitor.scala 629:69:chipyard.TestHarness.RocketConfig.fir@104757.4]
  wire [5:0] _T_1343; // @[Monitor.scala 629:69:chipyard.TestHarness.RocketConfig.fir@104757.4]
  wire [19:0] _T_1344; // @[Monitor.scala 629:44:chipyard.TestHarness.RocketConfig.fir@104758.4]
  wire [15:0] _T_1348; // @[Monitor.scala 606:57:chipyard.TestHarness.RocketConfig.fir@104762.4]
  wire [19:0] _GEN_74; // @[Monitor.scala 629:97:chipyard.TestHarness.RocketConfig.fir@104763.4]
  wire [19:0] _T_1349; // @[Monitor.scala 629:97:chipyard.TestHarness.RocketConfig.fir@104763.4]
  wire [19:0] _T_1350; // @[Monitor.scala 629:152:chipyard.TestHarness.RocketConfig.fir@104764.4]
  wire [19:0] _T_1352; // @[Monitor.scala 633:40:chipyard.TestHarness.RocketConfig.fir@104769.4]
  wire [19:0] _T_1357; // @[Monitor.scala 633:91:chipyard.TestHarness.RocketConfig.fir@104774.4]
  wire [19:0] _T_1358; // @[Monitor.scala 633:144:chipyard.TestHarness.RocketConfig.fir@104775.4]
  wire  _T_1362; // @[Monitor.scala 643:27:chipyard.TestHarness.RocketConfig.fir@104800.4]
  wire [7:0] _T_1364; // @[OneHot.scala 58:35:chipyard.TestHarness.RocketConfig.fir@104803.6]
  wire [3:0] _T_1365; // @[Monitor.scala 645:53:chipyard.TestHarness.RocketConfig.fir@104805.6]
  wire [3:0] _T_1366; // @[Monitor.scala 645:61:chipyard.TestHarness.RocketConfig.fir@104806.6]
  wire [3:0] _T_1367; // @[Monitor.scala 646:49:chipyard.TestHarness.RocketConfig.fir@104808.6]
  wire [3:0] _T_1368; // @[Monitor.scala 646:57:chipyard.TestHarness.RocketConfig.fir@104809.6]
  wire [4:0] _GEN_79; // @[Monitor.scala 647:72:chipyard.TestHarness.RocketConfig.fir@104811.6]
  wire [5:0] _T_1369; // @[Monitor.scala 647:72:chipyard.TestHarness.RocketConfig.fir@104811.6]
  wire [3:0] a_opcodes_set_interm; // @[Monitor.scala 643:72:chipyard.TestHarness.RocketConfig.fir@104802.4]
  wire [66:0] _GEN_80; // @[Monitor.scala 647:47:chipyard.TestHarness.RocketConfig.fir@104812.6]
  wire [66:0] _T_1370; // @[Monitor.scala 647:47:chipyard.TestHarness.RocketConfig.fir@104812.6]
  wire [3:0] a_sizes_set_interm; // @[Monitor.scala 643:72:chipyard.TestHarness.RocketConfig.fir@104802.4]
  wire [66:0] _GEN_82; // @[Monitor.scala 648:43:chipyard.TestHarness.RocketConfig.fir@104815.6]
  wire [66:0] _T_1372; // @[Monitor.scala 648:43:chipyard.TestHarness.RocketConfig.fir@104815.6]
  wire [4:0] _T_1373; // @[Monitor.scala 649:26:chipyard.TestHarness.RocketConfig.fir@104817.6]
  wire  _T_1375; // @[Monitor.scala 649:17:chipyard.TestHarness.RocketConfig.fir@104819.6]
  wire  _T_1377; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104821.6]
  wire  _T_1378; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104822.6]
  wire [7:0] _GEN_27; // @[Monitor.scala 643:72:chipyard.TestHarness.RocketConfig.fir@104802.4]
  wire [66:0] _GEN_30; // @[Monitor.scala 643:72:chipyard.TestHarness.RocketConfig.fir@104802.4]
  wire [66:0] _GEN_31; // @[Monitor.scala 643:72:chipyard.TestHarness.RocketConfig.fir@104802.4]
  wire  _T_1381; // @[Monitor.scala 660:27:chipyard.TestHarness.RocketConfig.fir@104836.4]
  wire  _T_1383; // @[Monitor.scala 660:75:chipyard.TestHarness.RocketConfig.fir@104838.4]
  wire  _T_1384; // @[Monitor.scala 660:72:chipyard.TestHarness.RocketConfig.fir@104839.4]
  wire [7:0] _T_1385; // @[OneHot.scala 58:35:chipyard.TestHarness.RocketConfig.fir@104841.6]
  wire [78:0] _GEN_84; // @[Monitor.scala 662:76:chipyard.TestHarness.RocketConfig.fir@104848.6]
  wire [78:0] _T_1391; // @[Monitor.scala 662:76:chipyard.TestHarness.RocketConfig.fir@104848.6]
  wire [7:0] _GEN_32; // @[Monitor.scala 660:91:chipyard.TestHarness.RocketConfig.fir@104840.4]
  wire [78:0] _GEN_33; // @[Monitor.scala 660:91:chipyard.TestHarness.RocketConfig.fir@104840.4]
  wire  _T_1398; // @[Monitor.scala 665:26:chipyard.TestHarness.RocketConfig.fir@104858.4]
  wire  _T_1401; // @[Monitor.scala 665:71:chipyard.TestHarness.RocketConfig.fir@104861.4]
  wire [4:0] _T_1402; // @[Monitor.scala 666:25:chipyard.TestHarness.RocketConfig.fir@104863.6]
  wire  _T_1404; // @[Monitor.scala 666:93:chipyard.TestHarness.RocketConfig.fir@104865.6]
  wire  _T_1405; // @[Monitor.scala 666:68:chipyard.TestHarness.RocketConfig.fir@104866.6]
  wire  _T_1406; // @[Monitor.scala 666:142:chipyard.TestHarness.RocketConfig.fir@104867.6]
  wire  _T_1407; // @[Monitor.scala 666:119:chipyard.TestHarness.RocketConfig.fir@104868.6]
  wire  _T_1408; // @[Monitor.scala 666:166:chipyard.TestHarness.RocketConfig.fir@104869.6]
  wire  _T_1409; // @[Monitor.scala 666:49:chipyard.TestHarness.RocketConfig.fir@104870.6]
  wire  _T_1411; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104872.6]
  wire  _T_1412; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104873.6]
  wire [3:0] a_opcode_lookup; // @[:chipyard.TestHarness.RocketConfig.fir@104755.4 :chipyard.TestHarness.RocketConfig.fir@104756.4 Monitor.scala 629:21:chipyard.TestHarness.RocketConfig.fir@104765.4]
  wire [2:0] _GEN_37; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  wire [2:0] _GEN_38; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  wire [2:0] _GEN_39; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  wire [2:0] _GEN_40; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  wire [2:0] _GEN_41; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  wire [2:0] _GEN_42; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  wire  _T_1414; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  wire [2:0] _GEN_49; // @[Monitor.scala 667:96:chipyard.TestHarness.RocketConfig.fir@104881.6]
  wire [2:0] _GEN_50; // @[Monitor.scala 667:96:chipyard.TestHarness.RocketConfig.fir@104881.6]
  wire  _T_1416; // @[Monitor.scala 667:96:chipyard.TestHarness.RocketConfig.fir@104881.6]
  wire  _T_1417; // @[Monitor.scala 667:71:chipyard.TestHarness.RocketConfig.fir@104882.6]
  wire [2:0] _GEN_53; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  wire [2:0] _GEN_54; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  wire [2:0] _GEN_55; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  wire [2:0] _GEN_56; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  wire [2:0] _GEN_57; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  wire [2:0] _GEN_58; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  wire  _T_1418; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  wire [2:0] _GEN_65; // @[Monitor.scala 668:124:chipyard.TestHarness.RocketConfig.fir@104884.6]
  wire [2:0] _GEN_66; // @[Monitor.scala 668:124:chipyard.TestHarness.RocketConfig.fir@104884.6]
  wire  _T_1419; // @[Monitor.scala 668:124:chipyard.TestHarness.RocketConfig.fir@104884.6]
  wire  _T_1420; // @[Monitor.scala 668:99:chipyard.TestHarness.RocketConfig.fir@104885.6]
  wire  _T_1421; // @[Monitor.scala 668:34:chipyard.TestHarness.RocketConfig.fir@104886.6]
  wire  _T_1422; // @[Monitor.scala 668:15:chipyard.TestHarness.RocketConfig.fir@104887.6]
  wire  _T_1424; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104889.6]
  wire  _T_1425; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104890.6]
  wire [3:0] a_size_lookup; // @[:chipyard.TestHarness.RocketConfig.fir@104766.4 :chipyard.TestHarness.RocketConfig.fir@104767.4 Monitor.scala 633:19:chipyard.TestHarness.RocketConfig.fir@104776.4]
  wire [3:0] _GEN_87; // @[Monitor.scala 670:34:chipyard.TestHarness.RocketConfig.fir@104895.6]
  wire  _T_1426; // @[Monitor.scala 670:34:chipyard.TestHarness.RocketConfig.fir@104895.6]
  wire  _T_1428; // @[Monitor.scala 670:72:chipyard.TestHarness.RocketConfig.fir@104897.6]
  wire  _T_1429; // @[Monitor.scala 670:53:chipyard.TestHarness.RocketConfig.fir@104898.6]
  wire  _T_1431; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104900.6]
  wire  _T_1432; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104901.6]
  wire  _T_1434; // @[Monitor.scala 672:36:chipyard.TestHarness.RocketConfig.fir@104908.4]
  wire  _T_1435; // @[Monitor.scala 672:47:chipyard.TestHarness.RocketConfig.fir@104909.4]
  wire  _T_1437; // @[Monitor.scala 672:65:chipyard.TestHarness.RocketConfig.fir@104911.4]
  wire  _T_1439; // @[Monitor.scala 672:116:chipyard.TestHarness.RocketConfig.fir@104913.4]
  wire  _T_1440; // @[Monitor.scala 673:15:chipyard.TestHarness.RocketConfig.fir@104915.6]
  wire  _T_1441; // @[Monitor.scala 673:32:chipyard.TestHarness.RocketConfig.fir@104916.6]
  wire  _T_1443; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104918.6]
  wire  _T_1444; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104919.6]
  wire [4:0] a_set; // @[:chipyard.TestHarness.RocketConfig.fir@104749.4 :chipyard.TestHarness.RocketConfig.fir@104750.4 Monitor.scala 644:13:chipyard.TestHarness.RocketConfig.fir@104804.6]
  wire [4:0] d_clr; // @[:chipyard.TestHarness.RocketConfig.fir@104828.4 :chipyard.TestHarness.RocketConfig.fir@104829.4 Monitor.scala 661:13:chipyard.TestHarness.RocketConfig.fir@104842.6]
  wire  _T_1445; // @[Monitor.scala 677:20:chipyard.TestHarness.RocketConfig.fir@104925.4]
  wire  _T_1446; // @[Monitor.scala 677:40:chipyard.TestHarness.RocketConfig.fir@104926.4]
  wire  _T_1447; // @[Monitor.scala 677:33:chipyard.TestHarness.RocketConfig.fir@104927.4]
  wire  _T_1448; // @[Monitor.scala 677:30:chipyard.TestHarness.RocketConfig.fir@104928.4]
  wire  _T_1450; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104930.4]
  wire  _T_1451; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104931.4]
  wire [4:0] _T_1452; // @[Monitor.scala 680:27:chipyard.TestHarness.RocketConfig.fir@104936.4]
  wire [4:0] _T_1453; // @[Monitor.scala 680:38:chipyard.TestHarness.RocketConfig.fir@104937.4]
  wire [4:0] _T_1454; // @[Monitor.scala 680:36:chipyard.TestHarness.RocketConfig.fir@104938.4]
  wire [19:0] a_opcodes_set; // @[:chipyard.TestHarness.RocketConfig.fir@104751.4 :chipyard.TestHarness.RocketConfig.fir@104752.4 Monitor.scala 647:21:chipyard.TestHarness.RocketConfig.fir@104813.6]
  wire [19:0] _T_1455; // @[Monitor.scala 681:43:chipyard.TestHarness.RocketConfig.fir@104940.4]
  wire [19:0] d_opcodes_clr; // @[:chipyard.TestHarness.RocketConfig.fir@104830.4 :chipyard.TestHarness.RocketConfig.fir@104831.4 Monitor.scala 662:21:chipyard.TestHarness.RocketConfig.fir@104849.6]
  wire [19:0] _T_1456; // @[Monitor.scala 681:62:chipyard.TestHarness.RocketConfig.fir@104941.4]
  wire [19:0] _T_1457; // @[Monitor.scala 681:60:chipyard.TestHarness.RocketConfig.fir@104942.4]
  wire [19:0] a_sizes_set; // @[:chipyard.TestHarness.RocketConfig.fir@104753.4 :chipyard.TestHarness.RocketConfig.fir@104754.4 Monitor.scala 648:19:chipyard.TestHarness.RocketConfig.fir@104816.6]
  wire [19:0] _T_1458; // @[Monitor.scala 682:39:chipyard.TestHarness.RocketConfig.fir@104944.4]
  wire [19:0] _T_1460; // @[Monitor.scala 682:54:chipyard.TestHarness.RocketConfig.fir@104946.4]
  reg [31:0] _T_1461; // @[Monitor.scala 684:27:chipyard.TestHarness.RocketConfig.fir@104948.4]
  reg [31:0] _RAND_27;
  wire  _T_1462; // @[Monitor.scala 687:26:chipyard.TestHarness.RocketConfig.fir@104951.4]
  wire  _T_1463; // @[Monitor.scala 687:16:chipyard.TestHarness.RocketConfig.fir@104952.4]
  wire  _T_1464; // @[Monitor.scala 687:39:chipyard.TestHarness.RocketConfig.fir@104953.4]
  wire  _T_1465; // @[Monitor.scala 687:30:chipyard.TestHarness.RocketConfig.fir@104954.4]
  wire  _T_1466; // @[Monitor.scala 687:59:chipyard.TestHarness.RocketConfig.fir@104955.4]
  wire  _T_1467; // @[Monitor.scala 687:47:chipyard.TestHarness.RocketConfig.fir@104956.4]
  wire  _T_1469; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104958.4]
  wire  _T_1470; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104959.4]
  wire [31:0] _T_1472; // @[Monitor.scala 689:26:chipyard.TestHarness.RocketConfig.fir@104965.4]
  wire  _T_1475; // @[Monitor.scala 690:27:chipyard.TestHarness.RocketConfig.fir@104969.4]
  reg [6:0] _T_1476; // @[Monitor.scala 694:27:chipyard.TestHarness.RocketConfig.fir@104973.4]
  reg [31:0] _RAND_28;
  reg [2:0] _T_1485; // @[Edges.scala 230:27:chipyard.TestHarness.RocketConfig.fir@104982.4]
  reg [31:0] _RAND_29;
  wire [2:0] _T_1487; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104984.4]
  wire  _T_1488; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104985.4]
  wire  _T_1498; // @[Monitor.scala 700:27:chipyard.TestHarness.RocketConfig.fir@104999.4]
  wire  _T_1501; // @[Edges.scala 72:43:chipyard.TestHarness.RocketConfig.fir@105002.4]
  wire  _T_1502; // @[Edges.scala 72:40:chipyard.TestHarness.RocketConfig.fir@105003.4]
  wire  _T_1503; // @[Monitor.scala 700:38:chipyard.TestHarness.RocketConfig.fir@105004.4]
  wire [7:0] _T_1504; // @[OneHot.scala 58:35:chipyard.TestHarness.RocketConfig.fir@105006.6]
  wire [6:0] _T_1505; // @[Monitor.scala 702:23:chipyard.TestHarness.RocketConfig.fir@105008.6]
  wire  _T_1507; // @[Monitor.scala 702:14:chipyard.TestHarness.RocketConfig.fir@105010.6]
  wire  _T_1509; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@105012.6]
  wire  _T_1510; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@105013.6]
  wire [7:0] _GEN_69; // @[Monitor.scala 700:72:chipyard.TestHarness.RocketConfig.fir@105005.4]
  wire [7:0] _T_1515; // @[OneHot.scala 58:35:chipyard.TestHarness.RocketConfig.fir@105025.6]
  wire [6:0] _T_1516; // @[Monitor.scala 708:24:chipyard.TestHarness.RocketConfig.fir@105027.6]
  wire [6:0] _T_1517; // @[Monitor.scala 708:35:chipyard.TestHarness.RocketConfig.fir@105028.6]
  wire  _T_1520; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@105031.6]
  wire  _T_1521; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@105032.6]
  wire [7:0] _GEN_70; // @[Monitor.scala 706:73:chipyard.TestHarness.RocketConfig.fir@105024.4]
  wire [6:0] _T_1522; // @[Monitor.scala 713:27:chipyard.TestHarness.RocketConfig.fir@105038.4]
  wire [6:0] _T_1523; // @[Monitor.scala 713:38:chipyard.TestHarness.RocketConfig.fir@105039.4]
  wire [6:0] _T_1524; // @[Monitor.scala 713:36:chipyard.TestHarness.RocketConfig.fir@105040.4]
  wire  _GEN_88; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102610.10]
  wire  _GEN_104; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102703.10]
  wire  _GEN_122; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102806.10]
  wire  _GEN_134; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102865.10]
  wire  _GEN_144; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102916.10]
  wire  _GEN_154; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102969.10]
  wire  _GEN_164; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103020.10]
  wire  _GEN_174; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103071.10]
  wire  _GEN_186; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103143.10]
  wire  _GEN_196; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103185.10]
  wire  _GEN_208; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103243.10]
  wire  _GEN_220; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103302.10]
  wire  _GEN_226; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103337.10]
  wire  _GEN_232; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103373.10]
  wire  _GEN_238; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104004.10]
  wire  _GEN_250; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104052.10]
  wire  _GEN_260; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104101.10]
  wire  _GEN_274; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104185.10]
  wire  _GEN_286; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104252.10]
  wire  _GEN_296; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104292.10]
  wire  _GEN_304; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104324.10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104949.4]
    .out(plusarg_reader_out)
  );
  assign _T_4 = io_in_a_bits_source == 3'h4; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@102470.6]
  assign _T_5 = io_in_a_bits_source == 3'h0; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@102471.6]
  assign _T_6 = io_in_a_bits_source == 3'h1; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@102472.6]
  assign _T_7 = io_in_a_bits_source == 3'h2; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@102473.6]
  assign _T_9 = _T_4 | _T_5; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@102480.6]
  assign _T_10 = _T_9 | _T_6; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@102481.6]
  assign _T_11 = _T_10 | _T_7; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@102482.6]
  assign _T_13 = 13'h3f << io_in_a_bits_size; // @[package.scala 189:77:chipyard.TestHarness.RocketConfig.fir@102484.6]
  assign _T_15 = ~_T_13[5:0]; // @[package.scala 189:46:chipyard.TestHarness.RocketConfig.fir@102486.6]
  assign _GEN_71 = {{26'd0}, _T_15}; // @[Edges.scala 22:16:chipyard.TestHarness.RocketConfig.fir@102487.6]
  assign _T_16 = io_in_a_bits_address & _GEN_71; // @[Edges.scala 22:16:chipyard.TestHarness.RocketConfig.fir@102487.6]
  assign _T_17 = _T_16 == 32'h0; // @[Edges.scala 22:24:chipyard.TestHarness.RocketConfig.fir@102488.6]
  assign _T_20 = 4'h1 << io_in_a_bits_size[1:0]; // @[OneHot.scala 65:12:chipyard.TestHarness.RocketConfig.fir@102491.6]
  assign _T_22 = _T_20[2:0] | 3'h1; // @[Misc.scala 201:81:chipyard.TestHarness.RocketConfig.fir@102493.6]
  assign _T_23 = io_in_a_bits_size >= 3'h3; // @[Misc.scala 205:21:chipyard.TestHarness.RocketConfig.fir@102494.6]
  assign _T_26 = ~io_in_a_bits_address[2]; // @[Misc.scala 210:20:chipyard.TestHarness.RocketConfig.fir@102497.6]
  assign _T_28 = _T_22[2] & _T_26; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102499.6]
  assign _T_29 = _T_23 | _T_28; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102500.6]
  assign _T_31 = _T_22[2] & io_in_a_bits_address[2]; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102502.6]
  assign _T_32 = _T_23 | _T_31; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102503.6]
  assign _T_35 = ~io_in_a_bits_address[1]; // @[Misc.scala 210:20:chipyard.TestHarness.RocketConfig.fir@102506.6]
  assign _T_36 = _T_26 & _T_35; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102507.6]
  assign _T_37 = _T_22[1] & _T_36; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102508.6]
  assign _T_38 = _T_29 | _T_37; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102509.6]
  assign _T_39 = _T_26 & io_in_a_bits_address[1]; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102510.6]
  assign _T_40 = _T_22[1] & _T_39; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102511.6]
  assign _T_41 = _T_29 | _T_40; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102512.6]
  assign _T_42 = io_in_a_bits_address[2] & _T_35; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102513.6]
  assign _T_43 = _T_22[1] & _T_42; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102514.6]
  assign _T_44 = _T_32 | _T_43; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102515.6]
  assign _T_45 = io_in_a_bits_address[2] & io_in_a_bits_address[1]; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102516.6]
  assign _T_46 = _T_22[1] & _T_45; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102517.6]
  assign _T_47 = _T_32 | _T_46; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102518.6]
  assign _T_50 = ~io_in_a_bits_address[0]; // @[Misc.scala 210:20:chipyard.TestHarness.RocketConfig.fir@102521.6]
  assign _T_51 = _T_36 & _T_50; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102522.6]
  assign _T_52 = _T_22[0] & _T_51; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102523.6]
  assign _T_53 = _T_38 | _T_52; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102524.6]
  assign _T_54 = _T_36 & io_in_a_bits_address[0]; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102525.6]
  assign _T_55 = _T_22[0] & _T_54; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102526.6]
  assign _T_56 = _T_38 | _T_55; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102527.6]
  assign _T_57 = _T_39 & _T_50; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102528.6]
  assign _T_58 = _T_22[0] & _T_57; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102529.6]
  assign _T_59 = _T_41 | _T_58; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102530.6]
  assign _T_60 = _T_39 & io_in_a_bits_address[0]; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102531.6]
  assign _T_61 = _T_22[0] & _T_60; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102532.6]
  assign _T_62 = _T_41 | _T_61; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102533.6]
  assign _T_63 = _T_42 & _T_50; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102534.6]
  assign _T_64 = _T_22[0] & _T_63; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102535.6]
  assign _T_65 = _T_44 | _T_64; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102536.6]
  assign _T_66 = _T_42 & io_in_a_bits_address[0]; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102537.6]
  assign _T_67 = _T_22[0] & _T_66; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102538.6]
  assign _T_68 = _T_44 | _T_67; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102539.6]
  assign _T_69 = _T_45 & _T_50; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102540.6]
  assign _T_70 = _T_22[0] & _T_69; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102541.6]
  assign _T_71 = _T_47 | _T_70; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102542.6]
  assign _T_72 = _T_45 & io_in_a_bits_address[0]; // @[Misc.scala 213:27:chipyard.TestHarness.RocketConfig.fir@102543.6]
  assign _T_73 = _T_22[0] & _T_72; // @[Misc.scala 214:38:chipyard.TestHarness.RocketConfig.fir@102544.6]
  assign _T_74 = _T_47 | _T_73; // @[Misc.scala 214:29:chipyard.TestHarness.RocketConfig.fir@102545.6]
  assign _T_81 = {_T_74,_T_71,_T_68,_T_65,_T_62,_T_59,_T_56,_T_53}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@102552.6]
  assign _T_120 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 79:25:chipyard.TestHarness.RocketConfig.fir@102595.6]
  assign _T_121 = 3'h6 == io_in_a_bits_size; // @[Parameters.scala 92:48:chipyard.TestHarness.RocketConfig.fir@102597.8]
  assign _T_123 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@102599.8]
  assign _T_124 = {1'b0,$signed(_T_123)}; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@102600.8]
  assign _T_126 = $signed(_T_124) & -33'sh10000000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@102602.8]
  assign _T_127 = $signed(_T_126) == 33'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@102603.8]
  assign _T_128 = _T_121 & _T_127; // @[Parameters.scala 551:56:chipyard.TestHarness.RocketConfig.fir@102604.8]
  assign _T_131 = _T_128 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102607.8]
  assign _T_132 = ~_T_131; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102608.8]
  assign _T_140 = _T_5 & _T_121; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@102625.8]
  assign _T_148 = _T_140 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102634.8]
  assign _T_149 = ~_T_148; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102635.8]
  assign _T_151 = _T_11 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102641.8]
  assign _T_152 = ~_T_151; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102642.8]
  assign _T_155 = _T_23 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102649.8]
  assign _T_156 = ~_T_155; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102650.8]
  assign _T_158 = _T_17 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102656.8]
  assign _T_159 = ~_T_158; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102657.8]
  assign _T_160 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 110:27:chipyard.TestHarness.RocketConfig.fir@102662.8]
  assign _T_162 = _T_160 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102664.8]
  assign _T_163 = ~_T_162; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102665.8]
  assign _T_164 = ~io_in_a_bits_mask; // @[Monitor.scala 86:18:chipyard.TestHarness.RocketConfig.fir@102670.8]
  assign _T_165 = _T_164 == 8'h0; // @[Monitor.scala 86:31:chipyard.TestHarness.RocketConfig.fir@102671.8]
  assign _T_167 = _T_165 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102673.8]
  assign _T_168 = ~_T_167; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102674.8]
  assign _T_169 = ~io_in_a_bits_corrupt; // @[Monitor.scala 87:18:chipyard.TestHarness.RocketConfig.fir@102679.8]
  assign _T_171 = _T_169 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102681.8]
  assign _T_172 = ~_T_171; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102682.8]
  assign _T_173 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 90:25:chipyard.TestHarness.RocketConfig.fir@102688.6]
  assign _T_217 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 97:31:chipyard.TestHarness.RocketConfig.fir@102763.8]
  assign _T_219 = _T_217 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102765.8]
  assign _T_220 = ~_T_219; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102766.8]
  assign _T_230 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 102:25:chipyard.TestHarness.RocketConfig.fir@102789.6]
  assign _T_232 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 93:42:chipyard.TestHarness.RocketConfig.fir@102792.8]
  assign _T_240 = _T_232 & _T_127; // @[Parameters.scala 551:56:chipyard.TestHarness.RocketConfig.fir@102800.8]
  assign _T_243 = _T_240 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102803.8]
  assign _T_244 = ~_T_243; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102804.8]
  assign _T_251 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 106:31:chipyard.TestHarness.RocketConfig.fir@102823.8]
  assign _T_253 = _T_251 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102825.8]
  assign _T_254 = ~_T_253; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102826.8]
  assign _T_255 = io_in_a_bits_mask == _T_81; // @[Monitor.scala 107:30:chipyard.TestHarness.RocketConfig.fir@102831.8]
  assign _T_257 = _T_255 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102833.8]
  assign _T_258 = ~_T_257; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102834.8]
  assign _T_263 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 111:25:chipyard.TestHarness.RocketConfig.fir@102848.6]
  assign _T_292 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 119:25:chipyard.TestHarness.RocketConfig.fir@102899.6]
  assign _T_317 = ~_T_81; // @[Monitor.scala 124:33:chipyard.TestHarness.RocketConfig.fir@102941.8]
  assign _T_318 = io_in_a_bits_mask & _T_317; // @[Monitor.scala 124:31:chipyard.TestHarness.RocketConfig.fir@102942.8]
  assign _T_319 = _T_318 == 8'h0; // @[Monitor.scala 124:40:chipyard.TestHarness.RocketConfig.fir@102943.8]
  assign _T_321 = _T_319 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102945.8]
  assign _T_322 = ~_T_321; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102946.8]
  assign _T_323 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 127:25:chipyard.TestHarness.RocketConfig.fir@102952.6]
  assign _T_325 = io_in_a_bits_size <= 3'h3; // @[Parameters.scala 93:42:chipyard.TestHarness.RocketConfig.fir@102955.8]
  assign _T_333 = _T_325 & _T_127; // @[Parameters.scala 551:56:chipyard.TestHarness.RocketConfig.fir@102963.8]
  assign _T_336 = _T_333 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102966.8]
  assign _T_337 = ~_T_336; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102967.8]
  assign _T_344 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 140:33:chipyard.TestHarness.RocketConfig.fir@102986.8]
  assign _T_346 = _T_344 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102988.8]
  assign _T_347 = ~_T_346; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102989.8]
  assign _T_352 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 135:25:chipyard.TestHarness.RocketConfig.fir@103003.6]
  assign _T_373 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 147:30:chipyard.TestHarness.RocketConfig.fir@103037.8]
  assign _T_375 = _T_373 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103039.8]
  assign _T_376 = ~_T_375; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103040.8]
  assign _T_381 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 143:25:chipyard.TestHarness.RocketConfig.fir@103054.6]
  assign _T_402 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 160:28:chipyard.TestHarness.RocketConfig.fir@103088.8]
  assign _T_404 = _T_402 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103090.8]
  assign _T_405 = ~_T_404; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103091.8]
  assign _T_414 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 44:24:chipyard.TestHarness.RocketConfig.fir@103115.6]
  assign _T_416 = _T_414 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103117.6]
  assign _T_417 = ~_T_416; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103118.6]
  assign _T_418 = io_in_d_bits_source == 3'h4; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103123.6]
  assign _T_419 = io_in_d_bits_source == 3'h0; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103124.6]
  assign _T_420 = io_in_d_bits_source == 3'h1; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103125.6]
  assign _T_421 = io_in_d_bits_source == 3'h2; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103126.6]
  assign _T_423 = _T_418 | _T_419; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@103133.6]
  assign _T_424 = _T_423 | _T_420; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@103134.6]
  assign _T_425 = _T_424 | _T_421; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@103135.6]
  assign _T_426 = io_in_d_bits_sink < 3'h7; // @[Monitor.scala 303:31:chipyard.TestHarness.RocketConfig.fir@103136.6]
  assign _T_427 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 307:25:chipyard.TestHarness.RocketConfig.fir@103137.6]
  assign _T_429 = _T_425 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103140.8]
  assign _T_430 = ~_T_429; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103141.8]
  assign _T_431 = io_in_d_bits_size >= 3'h3; // @[Monitor.scala 309:27:chipyard.TestHarness.RocketConfig.fir@103146.8]
  assign _T_433 = _T_431 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103148.8]
  assign _T_434 = ~_T_433; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103149.8]
  assign _T_435 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 310:28:chipyard.TestHarness.RocketConfig.fir@103154.8]
  assign _T_437 = _T_435 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103156.8]
  assign _T_438 = ~_T_437; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103157.8]
  assign _T_439 = ~io_in_d_bits_corrupt; // @[Monitor.scala 311:15:chipyard.TestHarness.RocketConfig.fir@103162.8]
  assign _T_441 = _T_439 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103164.8]
  assign _T_442 = ~_T_441; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103165.8]
  assign _T_443 = ~io_in_d_bits_denied; // @[Monitor.scala 312:15:chipyard.TestHarness.RocketConfig.fir@103170.8]
  assign _T_445 = _T_443 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103172.8]
  assign _T_446 = ~_T_445; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103173.8]
  assign _T_447 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 315:25:chipyard.TestHarness.RocketConfig.fir@103179.6]
  assign _T_452 = _T_426 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103189.8]
  assign _T_453 = ~_T_452; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103190.8]
  assign _T_458 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 104:26:chipyard.TestHarness.RocketConfig.fir@103203.8]
  assign _T_460 = _T_458 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103205.8]
  assign _T_461 = ~_T_460; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103206.8]
  assign _T_462 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 320:28:chipyard.TestHarness.RocketConfig.fir@103211.8]
  assign _T_464 = _T_462 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103213.8]
  assign _T_465 = ~_T_464; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103214.8]
  assign _T_475 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 325:25:chipyard.TestHarness.RocketConfig.fir@103237.6]
  assign _T_495 = _T_443 | io_in_d_bits_corrupt; // @[Monitor.scala 331:30:chipyard.TestHarness.RocketConfig.fir@103278.8]
  assign _T_497 = _T_495 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103280.8]
  assign _T_498 = ~_T_497; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103281.8]
  assign _T_504 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 335:25:chipyard.TestHarness.RocketConfig.fir@103296.6]
  assign _T_521 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 343:25:chipyard.TestHarness.RocketConfig.fir@103331.6]
  assign _T_539 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 351:25:chipyard.TestHarness.RocketConfig.fir@103367.6]
  assign _T_598 = io_in_b_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@103454.6]
  assign _T_599 = {1'b0,$signed(_T_598)}; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@103455.6]
  assign _T_601 = $signed(_T_599) & -33'sh10000000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@103457.6]
  assign _T_602 = $signed(_T_601) == 33'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@103458.6]
  assign _T_608 = io_in_b_bits_address & 32'h3f; // @[Edges.scala 22:16:chipyard.TestHarness.RocketConfig.fir@103466.6]
  assign _T_609 = _T_608 == 32'h0; // @[Edges.scala 22:24:chipyard.TestHarness.RocketConfig.fir@103467.6]
  assign _T_707 = _T_602 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103582.8]
  assign _T_708 = ~_T_707; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103583.8]
  assign _T_713 = _T_609 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103596.8]
  assign _T_714 = ~_T_713; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103597.8]
  assign _T_715 = io_in_b_bits_param <= 2'h2; // @[Bundles.scala 104:26:chipyard.TestHarness.RocketConfig.fir@103602.8]
  assign _T_717 = _T_715 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103604.8]
  assign _T_718 = ~_T_717; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103605.8]
  assign _T_863 = io_in_c_bits_source == 3'h4; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103929.6]
  assign _T_864 = io_in_c_bits_source == 3'h0; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103930.6]
  assign _T_865 = io_in_c_bits_source == 3'h1; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103931.6]
  assign _T_866 = io_in_c_bits_source == 3'h2; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@103932.6]
  assign _T_868 = _T_863 | _T_864; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@103939.6]
  assign _T_869 = _T_868 | _T_865; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@103940.6]
  assign _T_870 = _T_869 | _T_866; // @[Parameters.scala 924:46:chipyard.TestHarness.RocketConfig.fir@103941.6]
  assign _T_872 = 13'h3f << io_in_c_bits_size; // @[package.scala 189:77:chipyard.TestHarness.RocketConfig.fir@103943.6]
  assign _T_874 = ~_T_872[5:0]; // @[package.scala 189:46:chipyard.TestHarness.RocketConfig.fir@103945.6]
  assign _GEN_72 = {{26'd0}, _T_874}; // @[Edges.scala 22:16:chipyard.TestHarness.RocketConfig.fir@103946.6]
  assign _T_875 = io_in_c_bits_address & _GEN_72; // @[Edges.scala 22:16:chipyard.TestHarness.RocketConfig.fir@103946.6]
  assign _T_876 = _T_875 == 32'h0; // @[Edges.scala 22:24:chipyard.TestHarness.RocketConfig.fir@103947.6]
  assign _T_877 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:chipyard.TestHarness.RocketConfig.fir@103948.6]
  assign _T_878 = {1'b0,$signed(_T_877)}; // @[Parameters.scala 137:49:chipyard.TestHarness.RocketConfig.fir@103949.6]
  assign _T_880 = $signed(_T_878) & -33'sh10000000; // @[Parameters.scala 137:52:chipyard.TestHarness.RocketConfig.fir@103951.6]
  assign _T_881 = $signed(_T_880) == 33'sh0; // @[Parameters.scala 137:67:chipyard.TestHarness.RocketConfig.fir@103952.6]
  assign _T_921 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 239:25:chipyard.TestHarness.RocketConfig.fir@103998.6]
  assign _T_923 = _T_881 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104001.8]
  assign _T_924 = ~_T_923; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104002.8]
  assign _T_926 = _T_870 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104008.8]
  assign _T_927 = ~_T_926; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104009.8]
  assign _T_928 = io_in_c_bits_size >= 3'h3; // @[Monitor.scala 242:30:chipyard.TestHarness.RocketConfig.fir@104014.8]
  assign _T_930 = _T_928 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104016.8]
  assign _T_931 = ~_T_930; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104017.8]
  assign _T_933 = _T_876 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104023.8]
  assign _T_934 = ~_T_933; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104024.8]
  assign _T_935 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 122:29:chipyard.TestHarness.RocketConfig.fir@104029.8]
  assign _T_937 = _T_935 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104031.8]
  assign _T_938 = ~_T_937; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104032.8]
  assign _T_939 = ~io_in_c_bits_corrupt; // @[Monitor.scala 245:18:chipyard.TestHarness.RocketConfig.fir@104037.8]
  assign _T_941 = _T_939 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104039.8]
  assign _T_942 = ~_T_941; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104040.8]
  assign _T_943 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 248:25:chipyard.TestHarness.RocketConfig.fir@104046.6]
  assign _T_961 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 256:25:chipyard.TestHarness.RocketConfig.fir@104086.6]
  assign _T_962 = 3'h6 == io_in_c_bits_size; // @[Parameters.scala 92:48:chipyard.TestHarness.RocketConfig.fir@104088.8]
  assign _T_969 = _T_962 & _T_881; // @[Parameters.scala 551:56:chipyard.TestHarness.RocketConfig.fir@104095.8]
  assign _T_972 = _T_969 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104098.8]
  assign _T_973 = ~_T_972; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104099.8]
  assign _T_981 = _T_864 & _T_962; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@104116.8]
  assign _T_989 = _T_981 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104125.8]
  assign _T_990 = ~_T_989; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104126.8]
  assign _T_1001 = io_in_c_bits_param <= 3'h2; // @[Bundles.scala 116:29:chipyard.TestHarness.RocketConfig.fir@104153.8]
  assign _T_1003 = _T_1001 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104155.8]
  assign _T_1004 = ~_T_1003; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104156.8]
  assign _T_1009 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 266:25:chipyard.TestHarness.RocketConfig.fir@104170.6]
  assign _T_1053 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 275:25:chipyard.TestHarness.RocketConfig.fir@104246.6]
  assign _T_1063 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 279:31:chipyard.TestHarness.RocketConfig.fir@104269.8]
  assign _T_1065 = _T_1063 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104271.8]
  assign _T_1066 = ~_T_1065; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104272.8]
  assign _T_1071 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 283:25:chipyard.TestHarness.RocketConfig.fir@104286.6]
  assign _T_1085 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 290:25:chipyard.TestHarness.RocketConfig.fir@104318.6]
  assign _T_1103 = io_in_e_bits_sink < 3'h7; // @[Monitor.scala 361:31:chipyard.TestHarness.RocketConfig.fir@104360.6]
  assign _T_1105 = _T_1103 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104362.6]
  assign _T_1106 = ~_T_1105; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104363.6]
  assign _T_1107 = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37:chipyard.TestHarness.RocketConfig.fir@104369.4]
  assign _T_1114 = ~io_in_a_bits_opcode[2]; // @[Edges.scala 93:28:chipyard.TestHarness.RocketConfig.fir@104376.4]
  assign _T_1118 = _T_1116 - 3'h1; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104380.4]
  assign _T_1119 = _T_1116 == 3'h0; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104381.4]
  assign _T_1132 = ~_T_1119; // @[Monitor.scala 386:22:chipyard.TestHarness.RocketConfig.fir@104397.4]
  assign _T_1133 = io_in_a_valid & _T_1132; // @[Monitor.scala 386:19:chipyard.TestHarness.RocketConfig.fir@104398.4]
  assign _T_1134 = io_in_a_bits_opcode == _T_1127; // @[Monitor.scala 387:32:chipyard.TestHarness.RocketConfig.fir@104400.6]
  assign _T_1136 = _T_1134 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104402.6]
  assign _T_1137 = ~_T_1136; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104403.6]
  assign _T_1138 = io_in_a_bits_param == _T_1128; // @[Monitor.scala 388:32:chipyard.TestHarness.RocketConfig.fir@104408.6]
  assign _T_1140 = _T_1138 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104410.6]
  assign _T_1141 = ~_T_1140; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104411.6]
  assign _T_1142 = io_in_a_bits_size == _T_1129; // @[Monitor.scala 389:32:chipyard.TestHarness.RocketConfig.fir@104416.6]
  assign _T_1144 = _T_1142 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104418.6]
  assign _T_1145 = ~_T_1144; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104419.6]
  assign _T_1146 = io_in_a_bits_source == _T_1130; // @[Monitor.scala 390:32:chipyard.TestHarness.RocketConfig.fir@104424.6]
  assign _T_1148 = _T_1146 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104426.6]
  assign _T_1149 = ~_T_1148; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104427.6]
  assign _T_1150 = io_in_a_bits_address == _T_1131; // @[Monitor.scala 391:32:chipyard.TestHarness.RocketConfig.fir@104432.6]
  assign _T_1152 = _T_1150 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104434.6]
  assign _T_1153 = ~_T_1152; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104435.6]
  assign _T_1155 = _T_1107 & _T_1119; // @[Monitor.scala 393:20:chipyard.TestHarness.RocketConfig.fir@104442.4]
  assign _T_1156 = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37:chipyard.TestHarness.RocketConfig.fir@104450.4]
  assign _T_1158 = 13'h3f << io_in_d_bits_size; // @[package.scala 189:77:chipyard.TestHarness.RocketConfig.fir@104452.4]
  assign _T_1160 = ~_T_1158[5:0]; // @[package.scala 189:46:chipyard.TestHarness.RocketConfig.fir@104454.4]
  assign _T_1166 = _T_1164 - 3'h1; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104460.4]
  assign _T_1167 = _T_1164 == 3'h0; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104461.4]
  assign _T_1181 = ~_T_1167; // @[Monitor.scala 538:22:chipyard.TestHarness.RocketConfig.fir@104478.4]
  assign _T_1182 = io_in_d_valid & _T_1181; // @[Monitor.scala 538:19:chipyard.TestHarness.RocketConfig.fir@104479.4]
  assign _T_1183 = io_in_d_bits_opcode == _T_1175; // @[Monitor.scala 539:29:chipyard.TestHarness.RocketConfig.fir@104481.6]
  assign _T_1185 = _T_1183 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104483.6]
  assign _T_1186 = ~_T_1185; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104484.6]
  assign _T_1187 = io_in_d_bits_param == _T_1176; // @[Monitor.scala 540:29:chipyard.TestHarness.RocketConfig.fir@104489.6]
  assign _T_1189 = _T_1187 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104491.6]
  assign _T_1190 = ~_T_1189; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104492.6]
  assign _T_1191 = io_in_d_bits_size == _T_1177; // @[Monitor.scala 541:29:chipyard.TestHarness.RocketConfig.fir@104497.6]
  assign _T_1193 = _T_1191 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104499.6]
  assign _T_1194 = ~_T_1193; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104500.6]
  assign _T_1195 = io_in_d_bits_source == _T_1178; // @[Monitor.scala 542:29:chipyard.TestHarness.RocketConfig.fir@104505.6]
  assign _T_1197 = _T_1195 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104507.6]
  assign _T_1198 = ~_T_1197; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104508.6]
  assign _T_1199 = io_in_d_bits_sink == _T_1179; // @[Monitor.scala 543:29:chipyard.TestHarness.RocketConfig.fir@104513.6]
  assign _T_1201 = _T_1199 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104515.6]
  assign _T_1202 = ~_T_1201; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104516.6]
  assign _T_1203 = io_in_d_bits_denied == _T_1180; // @[Monitor.scala 544:29:chipyard.TestHarness.RocketConfig.fir@104521.6]
  assign _T_1205 = _T_1203 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104523.6]
  assign _T_1206 = ~_T_1205; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104524.6]
  assign _T_1208 = _T_1156 & _T_1167; // @[Monitor.scala 546:20:chipyard.TestHarness.RocketConfig.fir@104531.4]
  assign _T_1209 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37:chipyard.TestHarness.RocketConfig.fir@104540.4]
  assign _T_1220 = _T_1218 - 3'h1; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104551.4]
  assign _T_1221 = _T_1218 == 3'h0; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104552.4]
  assign _T_1234 = ~_T_1221; // @[Monitor.scala 409:22:chipyard.TestHarness.RocketConfig.fir@104568.4]
  assign _T_1235 = io_in_b_valid & _T_1234; // @[Monitor.scala 409:19:chipyard.TestHarness.RocketConfig.fir@104569.4]
  assign _T_1240 = io_in_b_bits_param == _T_1230; // @[Monitor.scala 411:32:chipyard.TestHarness.RocketConfig.fir@104579.6]
  assign _T_1242 = _T_1240 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104581.6]
  assign _T_1243 = ~_T_1242; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104582.6]
  assign _T_1252 = io_in_b_bits_address == _T_1233; // @[Monitor.scala 414:32:chipyard.TestHarness.RocketConfig.fir@104603.6]
  assign _T_1254 = _T_1252 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104605.6]
  assign _T_1255 = ~_T_1254; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104606.6]
  assign _T_1257 = _T_1209 & _T_1221; // @[Monitor.scala 416:20:chipyard.TestHarness.RocketConfig.fir@104613.4]
  assign _T_1258 = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37:chipyard.TestHarness.RocketConfig.fir@104621.4]
  assign _T_1268 = _T_1266 - 3'h1; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104631.4]
  assign _T_1269 = _T_1266 == 3'h0; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104632.4]
  assign _T_1282 = ~_T_1269; // @[Monitor.scala 514:22:chipyard.TestHarness.RocketConfig.fir@104648.4]
  assign _T_1283 = io_in_c_valid & _T_1282; // @[Monitor.scala 514:19:chipyard.TestHarness.RocketConfig.fir@104649.4]
  assign _T_1284 = io_in_c_bits_opcode == _T_1277; // @[Monitor.scala 515:32:chipyard.TestHarness.RocketConfig.fir@104651.6]
  assign _T_1286 = _T_1284 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104653.6]
  assign _T_1287 = ~_T_1286; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104654.6]
  assign _T_1288 = io_in_c_bits_param == _T_1278; // @[Monitor.scala 516:32:chipyard.TestHarness.RocketConfig.fir@104659.6]
  assign _T_1290 = _T_1288 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104661.6]
  assign _T_1291 = ~_T_1290; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104662.6]
  assign _T_1292 = io_in_c_bits_size == _T_1279; // @[Monitor.scala 517:32:chipyard.TestHarness.RocketConfig.fir@104667.6]
  assign _T_1294 = _T_1292 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104669.6]
  assign _T_1295 = ~_T_1294; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104670.6]
  assign _T_1296 = io_in_c_bits_source == _T_1280; // @[Monitor.scala 518:32:chipyard.TestHarness.RocketConfig.fir@104675.6]
  assign _T_1298 = _T_1296 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104677.6]
  assign _T_1299 = ~_T_1298; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104678.6]
  assign _T_1300 = io_in_c_bits_address == _T_1281; // @[Monitor.scala 519:32:chipyard.TestHarness.RocketConfig.fir@104683.6]
  assign _T_1302 = _T_1300 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104685.6]
  assign _T_1303 = ~_T_1302; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104686.6]
  assign _T_1305 = _T_1258 & _T_1269; // @[Monitor.scala 521:20:chipyard.TestHarness.RocketConfig.fir@104693.4]
  assign _T_1317 = _T_1315 - 3'h1; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104715.4]
  assign a_first = _T_1315 == 3'h0; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104716.4]
  assign _T_1335 = _T_1333 - 3'h1; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104737.4]
  assign d_first = _T_1333 == 3'h0; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104738.4]
  assign _GEN_73 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 629:69:chipyard.TestHarness.RocketConfig.fir@104757.4]
  assign _T_1343 = {{1'd0}, _GEN_73}; // @[Monitor.scala 629:69:chipyard.TestHarness.RocketConfig.fir@104757.4]
  assign _T_1344 = inflight_opcodes >> _T_1343; // @[Monitor.scala 629:44:chipyard.TestHarness.RocketConfig.fir@104758.4]
  assign _T_1348 = 16'h10 - 16'h1; // @[Monitor.scala 606:57:chipyard.TestHarness.RocketConfig.fir@104762.4]
  assign _GEN_74 = {{4'd0}, _T_1348}; // @[Monitor.scala 629:97:chipyard.TestHarness.RocketConfig.fir@104763.4]
  assign _T_1349 = _T_1344 & _GEN_74; // @[Monitor.scala 629:97:chipyard.TestHarness.RocketConfig.fir@104763.4]
  assign _T_1350 = {{1'd0}, _T_1349[19:1]}; // @[Monitor.scala 629:152:chipyard.TestHarness.RocketConfig.fir@104764.4]
  assign _T_1352 = inflight_sizes >> _T_1343; // @[Monitor.scala 633:40:chipyard.TestHarness.RocketConfig.fir@104769.4]
  assign _T_1357 = _T_1352 & _GEN_74; // @[Monitor.scala 633:91:chipyard.TestHarness.RocketConfig.fir@104774.4]
  assign _T_1358 = {{1'd0}, _T_1357[19:1]}; // @[Monitor.scala 633:144:chipyard.TestHarness.RocketConfig.fir@104775.4]
  assign _T_1362 = _T_1107 & a_first; // @[Monitor.scala 643:27:chipyard.TestHarness.RocketConfig.fir@104800.4]
  assign _T_1364 = 8'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35:chipyard.TestHarness.RocketConfig.fir@104803.6]
  assign _T_1365 = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 645:53:chipyard.TestHarness.RocketConfig.fir@104805.6]
  assign _T_1366 = _T_1365 | 4'h1; // @[Monitor.scala 645:61:chipyard.TestHarness.RocketConfig.fir@104806.6]
  assign _T_1367 = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 646:49:chipyard.TestHarness.RocketConfig.fir@104808.6]
  assign _T_1368 = _T_1367 | 4'h1; // @[Monitor.scala 646:57:chipyard.TestHarness.RocketConfig.fir@104809.6]
  assign _GEN_79 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 647:72:chipyard.TestHarness.RocketConfig.fir@104811.6]
  assign _T_1369 = {{1'd0}, _GEN_79}; // @[Monitor.scala 647:72:chipyard.TestHarness.RocketConfig.fir@104811.6]
  assign a_opcodes_set_interm = _T_1362 ? _T_1366 : 4'h0; // @[Monitor.scala 643:72:chipyard.TestHarness.RocketConfig.fir@104802.4]
  assign _GEN_80 = {{63'd0}, a_opcodes_set_interm}; // @[Monitor.scala 647:47:chipyard.TestHarness.RocketConfig.fir@104812.6]
  assign _T_1370 = _GEN_80 << _T_1369; // @[Monitor.scala 647:47:chipyard.TestHarness.RocketConfig.fir@104812.6]
  assign a_sizes_set_interm = _T_1362 ? _T_1368 : 4'h0; // @[Monitor.scala 643:72:chipyard.TestHarness.RocketConfig.fir@104802.4]
  assign _GEN_82 = {{63'd0}, a_sizes_set_interm}; // @[Monitor.scala 648:43:chipyard.TestHarness.RocketConfig.fir@104815.6]
  assign _T_1372 = _GEN_82 << _T_1369; // @[Monitor.scala 648:43:chipyard.TestHarness.RocketConfig.fir@104815.6]
  assign _T_1373 = inflight >> io_in_a_bits_source; // @[Monitor.scala 649:26:chipyard.TestHarness.RocketConfig.fir@104817.6]
  assign _T_1375 = ~_T_1373[0]; // @[Monitor.scala 649:17:chipyard.TestHarness.RocketConfig.fir@104819.6]
  assign _T_1377 = _T_1375 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104821.6]
  assign _T_1378 = ~_T_1377; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104822.6]
  assign _GEN_27 = _T_1362 ? _T_1364 : 8'h0; // @[Monitor.scala 643:72:chipyard.TestHarness.RocketConfig.fir@104802.4]
  assign _GEN_30 = _T_1362 ? _T_1370 : 67'h0; // @[Monitor.scala 643:72:chipyard.TestHarness.RocketConfig.fir@104802.4]
  assign _GEN_31 = _T_1362 ? _T_1372 : 67'h0; // @[Monitor.scala 643:72:chipyard.TestHarness.RocketConfig.fir@104802.4]
  assign _T_1381 = _T_1156 & d_first; // @[Monitor.scala 660:27:chipyard.TestHarness.RocketConfig.fir@104836.4]
  assign _T_1383 = ~_T_427; // @[Monitor.scala 660:75:chipyard.TestHarness.RocketConfig.fir@104838.4]
  assign _T_1384 = _T_1381 & _T_1383; // @[Monitor.scala 660:72:chipyard.TestHarness.RocketConfig.fir@104839.4]
  assign _T_1385 = 8'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35:chipyard.TestHarness.RocketConfig.fir@104841.6]
  assign _GEN_84 = {{63'd0}, _T_1348}; // @[Monitor.scala 662:76:chipyard.TestHarness.RocketConfig.fir@104848.6]
  assign _T_1391 = _GEN_84 << _T_1343; // @[Monitor.scala 662:76:chipyard.TestHarness.RocketConfig.fir@104848.6]
  assign _GEN_32 = _T_1384 ? _T_1385 : 8'h0; // @[Monitor.scala 660:91:chipyard.TestHarness.RocketConfig.fir@104840.4]
  assign _GEN_33 = _T_1384 ? _T_1391 : 79'h0; // @[Monitor.scala 660:91:chipyard.TestHarness.RocketConfig.fir@104840.4]
  assign _T_1398 = io_in_d_valid & d_first; // @[Monitor.scala 665:26:chipyard.TestHarness.RocketConfig.fir@104858.4]
  assign _T_1401 = _T_1398 & _T_1383; // @[Monitor.scala 665:71:chipyard.TestHarness.RocketConfig.fir@104861.4]
  assign _T_1402 = inflight >> io_in_d_bits_source; // @[Monitor.scala 666:25:chipyard.TestHarness.RocketConfig.fir@104863.6]
  assign _T_1404 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 666:93:chipyard.TestHarness.RocketConfig.fir@104865.6]
  assign _T_1405 = io_in_a_valid & _T_1404; // @[Monitor.scala 666:68:chipyard.TestHarness.RocketConfig.fir@104866.6]
  assign _T_1406 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 666:142:chipyard.TestHarness.RocketConfig.fir@104867.6]
  assign _T_1407 = _T_1405 & _T_1406; // @[Monitor.scala 666:119:chipyard.TestHarness.RocketConfig.fir@104868.6]
  assign _T_1408 = _T_1407 & a_first; // @[Monitor.scala 666:166:chipyard.TestHarness.RocketConfig.fir@104869.6]
  assign _T_1409 = _T_1402[0] | _T_1408; // @[Monitor.scala 666:49:chipyard.TestHarness.RocketConfig.fir@104870.6]
  assign _T_1411 = _T_1409 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104872.6]
  assign _T_1412 = ~_T_1411; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104873.6]
  assign a_opcode_lookup = _T_1350[3:0]; // @[:chipyard.TestHarness.RocketConfig.fir@104755.4 :chipyard.TestHarness.RocketConfig.fir@104756.4 Monitor.scala 629:21:chipyard.TestHarness.RocketConfig.fir@104765.4]
  assign _GEN_37 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  assign _GEN_38 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_37; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  assign _GEN_39 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_38; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  assign _GEN_40 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_39; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  assign _GEN_41 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_40; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  assign _GEN_42 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_41; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  assign _T_1414 = io_in_d_bits_opcode == _GEN_42; // @[Monitor.scala 667:37:chipyard.TestHarness.RocketConfig.fir@104879.6]
  assign _GEN_49 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_40; // @[Monitor.scala 667:96:chipyard.TestHarness.RocketConfig.fir@104881.6]
  assign _GEN_50 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_49; // @[Monitor.scala 667:96:chipyard.TestHarness.RocketConfig.fir@104881.6]
  assign _T_1416 = io_in_d_bits_opcode == _GEN_50; // @[Monitor.scala 667:96:chipyard.TestHarness.RocketConfig.fir@104881.6]
  assign _T_1417 = _T_1414 | _T_1416; // @[Monitor.scala 667:71:chipyard.TestHarness.RocketConfig.fir@104882.6]
  assign _GEN_53 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  assign _GEN_54 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_53; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  assign _GEN_55 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_54; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  assign _GEN_56 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_55; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  assign _GEN_57 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_56; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  assign _GEN_58 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_57; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  assign _T_1418 = io_in_d_bits_opcode == _GEN_58; // @[Monitor.scala 668:60:chipyard.TestHarness.RocketConfig.fir@104883.6]
  assign _GEN_65 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_56; // @[Monitor.scala 668:124:chipyard.TestHarness.RocketConfig.fir@104884.6]
  assign _GEN_66 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_65; // @[Monitor.scala 668:124:chipyard.TestHarness.RocketConfig.fir@104884.6]
  assign _T_1419 = io_in_d_bits_opcode == _GEN_66; // @[Monitor.scala 668:124:chipyard.TestHarness.RocketConfig.fir@104884.6]
  assign _T_1420 = _T_1418 | _T_1419; // @[Monitor.scala 668:99:chipyard.TestHarness.RocketConfig.fir@104885.6]
  assign _T_1421 = io_in_a_valid & _T_1420; // @[Monitor.scala 668:34:chipyard.TestHarness.RocketConfig.fir@104886.6]
  assign _T_1422 = _T_1417 | _T_1421; // @[Monitor.scala 668:15:chipyard.TestHarness.RocketConfig.fir@104887.6]
  assign _T_1424 = _T_1422 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104889.6]
  assign _T_1425 = ~_T_1424; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104890.6]
  assign a_size_lookup = _T_1358[3:0]; // @[:chipyard.TestHarness.RocketConfig.fir@104766.4 :chipyard.TestHarness.RocketConfig.fir@104767.4 Monitor.scala 633:19:chipyard.TestHarness.RocketConfig.fir@104776.4]
  assign _GEN_87 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 670:34:chipyard.TestHarness.RocketConfig.fir@104895.6]
  assign _T_1426 = _GEN_87 == a_size_lookup; // @[Monitor.scala 670:34:chipyard.TestHarness.RocketConfig.fir@104895.6]
  assign _T_1428 = io_in_a_valid & _T_1406; // @[Monitor.scala 670:72:chipyard.TestHarness.RocketConfig.fir@104897.6]
  assign _T_1429 = _T_1426 | _T_1428; // @[Monitor.scala 670:53:chipyard.TestHarness.RocketConfig.fir@104898.6]
  assign _T_1431 = _T_1429 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104900.6]
  assign _T_1432 = ~_T_1431; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104901.6]
  assign _T_1434 = _T_1398 & a_first; // @[Monitor.scala 672:36:chipyard.TestHarness.RocketConfig.fir@104908.4]
  assign _T_1435 = _T_1434 & io_in_a_valid; // @[Monitor.scala 672:47:chipyard.TestHarness.RocketConfig.fir@104909.4]
  assign _T_1437 = _T_1435 & _T_1404; // @[Monitor.scala 672:65:chipyard.TestHarness.RocketConfig.fir@104911.4]
  assign _T_1439 = _T_1437 & _T_1383; // @[Monitor.scala 672:116:chipyard.TestHarness.RocketConfig.fir@104913.4]
  assign _T_1440 = ~io_in_d_ready; // @[Monitor.scala 673:15:chipyard.TestHarness.RocketConfig.fir@104915.6]
  assign _T_1441 = _T_1440 | io_in_a_ready; // @[Monitor.scala 673:32:chipyard.TestHarness.RocketConfig.fir@104916.6]
  assign _T_1443 = _T_1441 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104918.6]
  assign _T_1444 = ~_T_1443; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104919.6]
  assign a_set = _GEN_27[4:0]; // @[:chipyard.TestHarness.RocketConfig.fir@104749.4 :chipyard.TestHarness.RocketConfig.fir@104750.4 Monitor.scala 644:13:chipyard.TestHarness.RocketConfig.fir@104804.6]
  assign d_clr = _GEN_32[4:0]; // @[:chipyard.TestHarness.RocketConfig.fir@104828.4 :chipyard.TestHarness.RocketConfig.fir@104829.4 Monitor.scala 661:13:chipyard.TestHarness.RocketConfig.fir@104842.6]
  assign _T_1445 = a_set != d_clr; // @[Monitor.scala 677:20:chipyard.TestHarness.RocketConfig.fir@104925.4]
  assign _T_1446 = |a_set; // @[Monitor.scala 677:40:chipyard.TestHarness.RocketConfig.fir@104926.4]
  assign _T_1447 = ~_T_1446; // @[Monitor.scala 677:33:chipyard.TestHarness.RocketConfig.fir@104927.4]
  assign _T_1448 = _T_1445 | _T_1447; // @[Monitor.scala 677:30:chipyard.TestHarness.RocketConfig.fir@104928.4]
  assign _T_1450 = _T_1448 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104930.4]
  assign _T_1451 = ~_T_1450; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104931.4]
  assign _T_1452 = inflight | a_set; // @[Monitor.scala 680:27:chipyard.TestHarness.RocketConfig.fir@104936.4]
  assign _T_1453 = ~d_clr; // @[Monitor.scala 680:38:chipyard.TestHarness.RocketConfig.fir@104937.4]
  assign _T_1454 = _T_1452 & _T_1453; // @[Monitor.scala 680:36:chipyard.TestHarness.RocketConfig.fir@104938.4]
  assign a_opcodes_set = _GEN_30[19:0]; // @[:chipyard.TestHarness.RocketConfig.fir@104751.4 :chipyard.TestHarness.RocketConfig.fir@104752.4 Monitor.scala 647:21:chipyard.TestHarness.RocketConfig.fir@104813.6]
  assign _T_1455 = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 681:43:chipyard.TestHarness.RocketConfig.fir@104940.4]
  assign d_opcodes_clr = _GEN_33[19:0]; // @[:chipyard.TestHarness.RocketConfig.fir@104830.4 :chipyard.TestHarness.RocketConfig.fir@104831.4 Monitor.scala 662:21:chipyard.TestHarness.RocketConfig.fir@104849.6]
  assign _T_1456 = ~d_opcodes_clr; // @[Monitor.scala 681:62:chipyard.TestHarness.RocketConfig.fir@104941.4]
  assign _T_1457 = _T_1455 & _T_1456; // @[Monitor.scala 681:60:chipyard.TestHarness.RocketConfig.fir@104942.4]
  assign a_sizes_set = _GEN_31[19:0]; // @[:chipyard.TestHarness.RocketConfig.fir@104753.4 :chipyard.TestHarness.RocketConfig.fir@104754.4 Monitor.scala 648:19:chipyard.TestHarness.RocketConfig.fir@104816.6]
  assign _T_1458 = inflight_sizes | a_sizes_set; // @[Monitor.scala 682:39:chipyard.TestHarness.RocketConfig.fir@104944.4]
  assign _T_1460 = _T_1458 & _T_1456; // @[Monitor.scala 682:54:chipyard.TestHarness.RocketConfig.fir@104946.4]
  assign _T_1462 = |inflight; // @[Monitor.scala 687:26:chipyard.TestHarness.RocketConfig.fir@104951.4]
  assign _T_1463 = ~_T_1462; // @[Monitor.scala 687:16:chipyard.TestHarness.RocketConfig.fir@104952.4]
  assign _T_1464 = plusarg_reader_out == 32'h0; // @[Monitor.scala 687:39:chipyard.TestHarness.RocketConfig.fir@104953.4]
  assign _T_1465 = _T_1463 | _T_1464; // @[Monitor.scala 687:30:chipyard.TestHarness.RocketConfig.fir@104954.4]
  assign _T_1466 = _T_1461 < plusarg_reader_out; // @[Monitor.scala 687:59:chipyard.TestHarness.RocketConfig.fir@104955.4]
  assign _T_1467 = _T_1465 | _T_1466; // @[Monitor.scala 687:47:chipyard.TestHarness.RocketConfig.fir@104956.4]
  assign _T_1469 = _T_1467 | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104958.4]
  assign _T_1470 = ~_T_1469; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104959.4]
  assign _T_1472 = _T_1461 + 32'h1; // @[Monitor.scala 689:26:chipyard.TestHarness.RocketConfig.fir@104965.4]
  assign _T_1475 = _T_1107 | _T_1156; // @[Monitor.scala 690:27:chipyard.TestHarness.RocketConfig.fir@104969.4]
  assign _T_1487 = _T_1485 - 3'h1; // @[Edges.scala 231:28:chipyard.TestHarness.RocketConfig.fir@104984.4]
  assign _T_1488 = _T_1485 == 3'h0; // @[Edges.scala 232:25:chipyard.TestHarness.RocketConfig.fir@104985.4]
  assign _T_1498 = _T_1156 & _T_1488; // @[Monitor.scala 700:27:chipyard.TestHarness.RocketConfig.fir@104999.4]
  assign _T_1501 = ~io_in_d_bits_opcode[1]; // @[Edges.scala 72:43:chipyard.TestHarness.RocketConfig.fir@105002.4]
  assign _T_1502 = io_in_d_bits_opcode[2] & _T_1501; // @[Edges.scala 72:40:chipyard.TestHarness.RocketConfig.fir@105003.4]
  assign _T_1503 = _T_1498 & _T_1502; // @[Monitor.scala 700:38:chipyard.TestHarness.RocketConfig.fir@105004.4]
  assign _T_1504 = 8'h1 << io_in_d_bits_sink; // @[OneHot.scala 58:35:chipyard.TestHarness.RocketConfig.fir@105006.6]
  assign _T_1505 = _T_1476 >> io_in_d_bits_sink; // @[Monitor.scala 702:23:chipyard.TestHarness.RocketConfig.fir@105008.6]
  assign _T_1507 = ~_T_1505[0]; // @[Monitor.scala 702:14:chipyard.TestHarness.RocketConfig.fir@105010.6]
  assign _T_1509 = _T_1507 | reset; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@105012.6]
  assign _T_1510 = ~_T_1509; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@105013.6]
  assign _GEN_69 = _T_1503 ? _T_1504 : 8'h0; // @[Monitor.scala 700:72:chipyard.TestHarness.RocketConfig.fir@105005.4]
  assign _T_1515 = 8'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35:chipyard.TestHarness.RocketConfig.fir@105025.6]
  assign _T_1516 = _GEN_69[6:0] | _T_1476; // @[Monitor.scala 708:24:chipyard.TestHarness.RocketConfig.fir@105027.6]
  assign _T_1517 = _T_1516 >> io_in_e_bits_sink; // @[Monitor.scala 708:35:chipyard.TestHarness.RocketConfig.fir@105028.6]
  assign _T_1520 = _T_1517[0] | reset; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@105031.6]
  assign _T_1521 = ~_T_1520; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@105032.6]
  assign _GEN_70 = io_in_e_valid ? _T_1515 : 8'h0; // @[Monitor.scala 706:73:chipyard.TestHarness.RocketConfig.fir@105024.4]
  assign _T_1522 = _T_1476 | _GEN_69[6:0]; // @[Monitor.scala 713:27:chipyard.TestHarness.RocketConfig.fir@105038.4]
  assign _T_1523 = ~_GEN_70[6:0]; // @[Monitor.scala 713:38:chipyard.TestHarness.RocketConfig.fir@105039.4]
  assign _T_1524 = _T_1522 & _T_1523; // @[Monitor.scala 713:36:chipyard.TestHarness.RocketConfig.fir@105040.4]
  assign _GEN_88 = io_in_a_valid & _T_120; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102610.10]
  assign _GEN_104 = io_in_a_valid & _T_173; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102703.10]
  assign _GEN_122 = io_in_a_valid & _T_230; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102806.10]
  assign _GEN_134 = io_in_a_valid & _T_263; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102865.10]
  assign _GEN_144 = io_in_a_valid & _T_292; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102916.10]
  assign _GEN_154 = io_in_a_valid & _T_323; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102969.10]
  assign _GEN_164 = io_in_a_valid & _T_352; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103020.10]
  assign _GEN_174 = io_in_a_valid & _T_381; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103071.10]
  assign _GEN_186 = io_in_d_valid & _T_427; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103143.10]
  assign _GEN_196 = io_in_d_valid & _T_447; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103185.10]
  assign _GEN_208 = io_in_d_valid & _T_475; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103243.10]
  assign _GEN_220 = io_in_d_valid & _T_504; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103302.10]
  assign _GEN_226 = io_in_d_valid & _T_521; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103337.10]
  assign _GEN_232 = io_in_d_valid & _T_539; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103373.10]
  assign _GEN_238 = io_in_c_valid & _T_921; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104004.10]
  assign _GEN_250 = io_in_c_valid & _T_943; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104052.10]
  assign _GEN_260 = io_in_c_valid & _T_961; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104101.10]
  assign _GEN_274 = io_in_c_valid & _T_1009; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104185.10]
  assign _GEN_286 = io_in_c_valid & _T_1053; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104252.10]
  assign _GEN_296 = io_in_c_valid & _T_1071; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104292.10]
  assign _GEN_304 = io_in_c_valid & _T_1085; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104324.10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1116 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1127 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1128 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1129 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1130 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1131 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1164 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1175 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1176 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1177 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1178 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_1179 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1180 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_1218 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_1230 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_1233 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1266 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_1277 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_1278 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_1279 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_1280 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_1281 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  inflight = _RAND_22[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  inflight_opcodes = _RAND_23[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  inflight_sizes = _RAND_24[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_1315 = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_1333 = _RAND_26[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_1461 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_1476 = _RAND_28[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_1485 = _RAND_29[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1116 <= 3'h0;
    end else if (_T_1107) begin
      if (_T_1119) begin
        if (_T_1114) begin
          _T_1116 <= _T_15[5:3];
        end else begin
          _T_1116 <= 3'h0;
        end
      end else begin
        _T_1116 <= _T_1118;
      end
    end
    if (_T_1155) begin
      _T_1127 <= io_in_a_bits_opcode;
    end
    if (_T_1155) begin
      _T_1128 <= io_in_a_bits_param;
    end
    if (_T_1155) begin
      _T_1129 <= io_in_a_bits_size;
    end
    if (_T_1155) begin
      _T_1130 <= io_in_a_bits_source;
    end
    if (_T_1155) begin
      _T_1131 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_1164 <= 3'h0;
    end else if (_T_1156) begin
      if (_T_1167) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1164 <= _T_1160[5:3];
        end else begin
          _T_1164 <= 3'h0;
        end
      end else begin
        _T_1164 <= _T_1166;
      end
    end
    if (_T_1208) begin
      _T_1175 <= io_in_d_bits_opcode;
    end
    if (_T_1208) begin
      _T_1176 <= io_in_d_bits_param;
    end
    if (_T_1208) begin
      _T_1177 <= io_in_d_bits_size;
    end
    if (_T_1208) begin
      _T_1178 <= io_in_d_bits_source;
    end
    if (_T_1208) begin
      _T_1179 <= io_in_d_bits_sink;
    end
    if (_T_1208) begin
      _T_1180 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_1218 <= 3'h0;
    end else if (_T_1209) begin
      if (_T_1221) begin
        _T_1218 <= 3'h0;
      end else begin
        _T_1218 <= _T_1220;
      end
    end
    if (_T_1257) begin
      _T_1230 <= io_in_b_bits_param;
    end
    if (_T_1257) begin
      _T_1233 <= io_in_b_bits_address;
    end
    if (reset) begin
      _T_1266 <= 3'h0;
    end else if (_T_1258) begin
      if (_T_1269) begin
        if (io_in_c_bits_opcode[0]) begin
          _T_1266 <= _T_874[5:3];
        end else begin
          _T_1266 <= 3'h0;
        end
      end else begin
        _T_1266 <= _T_1268;
      end
    end
    if (_T_1305) begin
      _T_1277 <= io_in_c_bits_opcode;
    end
    if (_T_1305) begin
      _T_1278 <= io_in_c_bits_param;
    end
    if (_T_1305) begin
      _T_1279 <= io_in_c_bits_size;
    end
    if (_T_1305) begin
      _T_1280 <= io_in_c_bits_source;
    end
    if (_T_1305) begin
      _T_1281 <= io_in_c_bits_address;
    end
    if (reset) begin
      inflight <= 5'h0;
    end else begin
      inflight <= _T_1454;
    end
    if (reset) begin
      inflight_opcodes <= 20'h0;
    end else begin
      inflight_opcodes <= _T_1457;
    end
    if (reset) begin
      inflight_sizes <= 20'h0;
    end else begin
      inflight_sizes <= _T_1460;
    end
    if (reset) begin
      _T_1315 <= 3'h0;
    end else if (_T_1107) begin
      if (a_first) begin
        if (_T_1114) begin
          _T_1315 <= _T_15[5:3];
        end else begin
          _T_1315 <= 3'h0;
        end
      end else begin
        _T_1315 <= _T_1317;
      end
    end
    if (reset) begin
      _T_1333 <= 3'h0;
    end else if (_T_1156) begin
      if (d_first) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1333 <= _T_1160[5:3];
        end else begin
          _T_1333 <= 3'h0;
        end
      end else begin
        _T_1333 <= _T_1335;
      end
    end
    if (reset) begin
      _T_1461 <= 32'h0;
    end else if (_T_1475) begin
      _T_1461 <= 32'h0;
    end else begin
      _T_1461 <= _T_1472;
    end
    if (reset) begin
      _T_1476 <= 7'h0;
    end else begin
      _T_1476 <= _T_1524;
    end
    if (reset) begin
      _T_1485 <= 3'h0;
    end else if (_T_1156) begin
      if (_T_1488) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1485 <= _T_1160[5:3];
        end else begin
          _T_1485 <= 3'h0;
        end
      end else begin
        _T_1485 <= _T_1487;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_88 & _T_132) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102610.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_88 & _T_132) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102611.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_88 & _T_149) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102637.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_88 & _T_149) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102638.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_88 & _T_152) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102644.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_88 & _T_152) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102645.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_88 & _T_156) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102652.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_88 & _T_156) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102653.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_88 & _T_159) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102659.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_88 & _T_159) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102660.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_88 & _T_163) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102667.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_88 & _T_163) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102668.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_88 & _T_168) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102676.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_88 & _T_168) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102677.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_88 & _T_172) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102684.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_88 & _T_172) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102685.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_104 & _T_132) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102703.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_104 & _T_132) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102704.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_104 & _T_149) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102730.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_104 & _T_149) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102731.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_104 & _T_152) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102737.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_104 & _T_152) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102738.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_104 & _T_156) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102745.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_104 & _T_156) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102746.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_104 & _T_159) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102752.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_104 & _T_159) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102753.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_104 & _T_163) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102760.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_104 & _T_163) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102761.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_104 & _T_220) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102768.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_104 & _T_220) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102769.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_104 & _T_168) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102777.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_104 & _T_168) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102778.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_104 & _T_172) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102785.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_104 & _T_172) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102786.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_244) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102806.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & _T_244) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102807.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_152) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102813.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & _T_152) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102814.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_159) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102820.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & _T_159) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102821.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_254) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102828.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & _T_254) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102829.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_258) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102836.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & _T_258) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102837.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_172) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102844.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & _T_172) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102845.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & _T_244) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102865.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & _T_244) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102866.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & _T_152) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102872.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & _T_152) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102873.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & _T_159) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102879.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & _T_159) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102880.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & _T_254) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102887.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & _T_254) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102888.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & _T_258) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102895.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & _T_258) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102896.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_244) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102916.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_244) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102917.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_152) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102923.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_152) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102924.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_159) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102930.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_159) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102931.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_254) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102938.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_254) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102939.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_322) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102948.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_322) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102949.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_154 & _T_337) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102969.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_154 & _T_337) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102970.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_154 & _T_152) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102976.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_154 & _T_152) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102977.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_154 & _T_159) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102983.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_154 & _T_159) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102984.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_154 & _T_347) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102991.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_154 & _T_347) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102992.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_154 & _T_258) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@102999.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_154 & _T_258) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103000.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_164 & _T_337) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103020.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_164 & _T_337) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103021.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_164 & _T_152) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103027.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_164 & _T_152) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103028.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_164 & _T_159) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103034.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_164 & _T_159) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103035.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_164 & _T_376) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103042.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_164 & _T_376) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103043.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_164 & _T_258) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103050.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_164 & _T_258) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103051.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_174 & _T_244) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103071.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_174 & _T_244) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103072.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_174 & _T_152) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103078.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_174 & _T_152) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103079.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_174 & _T_159) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103085.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_174 & _T_159) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103086.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_174 & _T_405) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid opcode param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103093.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_174 & _T_405) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103094.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_174 & _T_258) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103101.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_174 & _T_258) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103102.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_174 & _T_172) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103109.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_174 & _T_172) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103110.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_417) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103120.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_417) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103121.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_430) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103143.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_430) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103144.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_434) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103151.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_434) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103152.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_438) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103159.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_438) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103160.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_442) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103167.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_442) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103168.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_446) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103175.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_446) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103176.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_196 & _T_430) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103185.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_196 & _T_430) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103186.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_196 & _T_453) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103192.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_196 & _T_453) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103193.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_196 & _T_434) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103200.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_196 & _T_434) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103201.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_196 & _T_461) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103208.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_196 & _T_461) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103209.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_196 & _T_465) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103216.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_196 & _T_465) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103217.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_196 & _T_442) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103224.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_196 & _T_442) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103225.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_430) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103243.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_430) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103244.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_453) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103250.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_453) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103251.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_434) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103258.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_434) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103259.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_461) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103266.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_461) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103267.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_465) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103274.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_465) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103275.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_498) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103283.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_498) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103284.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_220 & _T_430) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103302.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_220 & _T_430) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103303.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_220 & _T_438) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103310.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_220 & _T_438) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103311.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_220 & _T_442) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103318.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_220 & _T_442) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103319.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_226 & _T_430) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103337.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_226 & _T_430) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103338.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_226 & _T_438) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103345.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_226 & _T_438) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103346.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_226 & _T_498) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103354.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_226 & _T_498) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103355.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_232 & _T_430) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103373.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_232 & _T_430) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103374.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_232 & _T_438) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103381.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_232 & _T_438) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103382.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_232 & _T_442) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103389.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_232 & _T_442) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@103390.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & _T_708) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103585.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & _T_708) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103586.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & _T_714) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103599.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & _T_714) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103600.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & _T_718) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103607.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & _T_718) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@103608.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_238 & _T_924) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104004.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_238 & _T_924) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104005.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_238 & _T_927) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104011.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_238 & _T_927) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104012.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_238 & _T_931) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104019.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_238 & _T_931) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104020.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_238 & _T_934) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104026.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_238 & _T_934) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104027.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_238 & _T_938) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104034.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_238 & _T_938) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104035.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_238 & _T_942) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck is corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104042.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_238 & _T_942) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104043.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_250 & _T_924) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104052.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_250 & _T_924) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104053.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_250 & _T_927) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104059.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_250 & _T_927) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104060.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_250 & _T_931) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104067.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_250 & _T_931) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104068.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_250 & _T_934) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104074.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_250 & _T_934) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104075.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_250 & _T_938) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104082.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_250 & _T_938) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104083.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_973) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104101.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_973) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104102.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_990) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104128.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_990) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104129.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_927) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104135.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_927) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104136.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_931) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104143.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_931) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104144.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_934) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104150.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_934) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104151.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_1004) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104158.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_1004) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104159.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_942) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release is corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104166.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_942) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104167.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_274 & _T_973) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104185.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_274 & _T_973) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104186.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_274 & _T_990) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104212.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_274 & _T_990) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104213.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_274 & _T_927) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104219.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_274 & _T_927) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104220.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_274 & _T_931) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104227.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_274 & _T_931) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104228.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_274 & _T_934) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104234.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_274 & _T_934) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104235.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_274 & _T_1004) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104242.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_274 & _T_1004) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104243.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_286 & _T_924) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104252.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_286 & _T_924) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104253.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_286 & _T_927) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104259.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_286 & _T_927) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104260.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_286 & _T_934) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104266.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_286 & _T_934) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104267.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_286 & _T_1066) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104274.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_286 & _T_1066) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104275.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_286 & _T_942) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck is corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104282.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_286 & _T_942) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104283.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_296 & _T_924) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104292.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_296 & _T_924) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104293.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_296 & _T_927) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104299.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_296 & _T_927) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104300.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_296 & _T_934) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104306.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_296 & _T_934) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104307.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_296 & _T_1066) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104314.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_296 & _T_1066) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104315.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_304 & _T_924) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104324.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_304 & _T_924) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104325.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_304 & _T_927) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104331.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_304 & _T_927) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104332.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_304 & _T_934) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104338.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_304 & _T_934) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104339.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_304 & _T_1066) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104346.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_304 & _T_1066) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104347.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_304 & _T_942) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck is corrupt (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104354.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_304 & _T_942) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104355.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & _T_1106) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channels carries invalid sink ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104365.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & _T_1106) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104366.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1133 & _T_1137) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104405.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1133 & _T_1137) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104406.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1133 & _T_1141) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104413.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1133 & _T_1141) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104414.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1133 & _T_1145) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104421.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1133 & _T_1145) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104422.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1133 & _T_1149) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104429.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1133 & _T_1149) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104430.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1133 & _T_1153) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104437.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1133 & _T_1153) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104438.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1182 & _T_1186) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104486.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1182 & _T_1186) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104487.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1182 & _T_1190) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104494.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1182 & _T_1190) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104495.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1182 & _T_1194) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104502.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1182 & _T_1194) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104503.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1182 & _T_1198) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104510.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1182 & _T_1198) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104511.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1182 & _T_1202) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104518.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1182 & _T_1202) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104519.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1182 & _T_1206) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104526.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1182 & _T_1206) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104527.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1235 & _T_1243) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104584.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1235 & _T_1243) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104585.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1235 & _T_1255) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104608.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1235 & _T_1255) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104609.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1283 & _T_1287) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104656.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1283 & _T_1287) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104657.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1283 & _T_1291) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104664.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1283 & _T_1291) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104665.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1283 & _T_1295) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104672.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1283 & _T_1295) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104673.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1283 & _T_1299) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104680.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1283 & _T_1299) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104681.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1283 & _T_1303) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104688.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1283 & _T_1303) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104689.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1362 & _T_1378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104824.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1362 & _T_1378) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104825.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1401 & _T_1412) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104875.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1401 & _T_1412) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104876.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1401 & _T_1425) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104892.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1401 & _T_1425) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104893.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1401 & _T_1432) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104903.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1401 & _T_1432) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104904.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1439 & _T_1444) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104921.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1439 & _T_1444) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104922.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1451) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 2 (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104933.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1451) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@104934.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1470) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104961.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1470) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@104962.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1510) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@105015.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1510) begin
          $fatal; // @[Monitor.scala 51:11:chipyard.TestHarness.RocketConfig.fir@105016.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & _T_1521) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at BankedL2Params.scala:58:27)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@105034.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & _T_1521) begin
          $fatal; // @[Monitor.scala 44:11:chipyard.TestHarness.RocketConfig.fir@105035.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
