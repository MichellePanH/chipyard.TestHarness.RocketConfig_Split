module INToRecFN( // @[:chipyard.TestHarness.RocketConfig.fir@235416.2]
  input         io_signedIn, // @[:chipyard.TestHarness.RocketConfig.fir@235417.4]
  input  [63:0] io_in, // @[:chipyard.TestHarness.RocketConfig.fir@235417.4]
  input  [2:0]  io_roundingMode, // @[:chipyard.TestHarness.RocketConfig.fir@235417.4]
  output [32:0] io_out, // @[:chipyard.TestHarness.RocketConfig.fir@235417.4]
  output [4:0]  io_exceptionFlags // @[:chipyard.TestHarness.RocketConfig.fir@235417.4]
);
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[INToRecFN.scala 59:15:chipyard.TestHarness.RocketConfig.fir@235570.4]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[INToRecFN.scala 59:15:chipyard.TestHarness.RocketConfig.fir@235570.4]
  wire [8:0] roundAnyRawFNToRecFN_io_in_sExp; // @[INToRecFN.scala 59:15:chipyard.TestHarness.RocketConfig.fir@235570.4]
  wire [64:0] roundAnyRawFNToRecFN_io_in_sig; // @[INToRecFN.scala 59:15:chipyard.TestHarness.RocketConfig.fir@235570.4]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[INToRecFN.scala 59:15:chipyard.TestHarness.RocketConfig.fir@235570.4]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 59:15:chipyard.TestHarness.RocketConfig.fir@235570.4]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 59:15:chipyard.TestHarness.RocketConfig.fir@235570.4]
  wire  intAsRawFloat_sign; // @[rawFloatFromIN.scala 50:29:chipyard.TestHarness.RocketConfig.fir@235421.4]
  wire [63:0] _T_3; // @[rawFloatFromIN.scala 51:31:chipyard.TestHarness.RocketConfig.fir@235423.4]
  wire [63:0] _T_4; // @[rawFloatFromIN.scala 51:24:chipyard.TestHarness.RocketConfig.fir@235424.4]
  wire [127:0] _T_5; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@235425.4]
  wire [5:0] _T_71; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235491.4]
  wire [5:0] _T_72; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235492.4]
  wire [5:0] _T_73; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235493.4]
  wire [5:0] _T_74; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235494.4]
  wire [5:0] _T_75; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235495.4]
  wire [5:0] _T_76; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235496.4]
  wire [5:0] _T_77; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235497.4]
  wire [5:0] _T_78; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235498.4]
  wire [5:0] _T_79; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235499.4]
  wire [5:0] _T_80; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235500.4]
  wire [5:0] _T_81; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235501.4]
  wire [5:0] _T_82; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235502.4]
  wire [5:0] _T_83; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235503.4]
  wire [5:0] _T_84; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235504.4]
  wire [5:0] _T_85; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235505.4]
  wire [5:0] _T_86; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235506.4]
  wire [5:0] _T_87; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235507.4]
  wire [5:0] _T_88; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235508.4]
  wire [5:0] _T_89; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235509.4]
  wire [5:0] _T_90; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235510.4]
  wire [5:0] _T_91; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235511.4]
  wire [5:0] _T_92; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235512.4]
  wire [5:0] _T_93; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235513.4]
  wire [5:0] _T_94; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235514.4]
  wire [5:0] _T_95; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235515.4]
  wire [5:0] _T_96; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235516.4]
  wire [5:0] _T_97; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235517.4]
  wire [5:0] _T_98; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235518.4]
  wire [5:0] _T_99; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235519.4]
  wire [5:0] _T_100; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235520.4]
  wire [5:0] _T_101; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235521.4]
  wire [5:0] _T_102; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235522.4]
  wire [5:0] _T_103; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235523.4]
  wire [5:0] _T_104; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235524.4]
  wire [5:0] _T_105; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235525.4]
  wire [5:0] _T_106; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235526.4]
  wire [5:0] _T_107; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235527.4]
  wire [5:0] _T_108; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235528.4]
  wire [5:0] _T_109; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235529.4]
  wire [5:0] _T_110; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235530.4]
  wire [5:0] _T_111; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235531.4]
  wire [5:0] _T_112; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235532.4]
  wire [5:0] _T_113; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235533.4]
  wire [5:0] _T_114; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235534.4]
  wire [5:0] _T_115; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235535.4]
  wire [5:0] _T_116; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235536.4]
  wire [5:0] _T_117; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235537.4]
  wire [5:0] _T_118; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235538.4]
  wire [5:0] _T_119; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235539.4]
  wire [5:0] _T_120; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235540.4]
  wire [5:0] _T_121; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235541.4]
  wire [5:0] _T_122; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235542.4]
  wire [5:0] _T_123; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235543.4]
  wire [5:0] _T_124; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235544.4]
  wire [5:0] _T_125; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235545.4]
  wire [5:0] _T_126; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235546.4]
  wire [5:0] _T_127; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235547.4]
  wire [5:0] _T_128; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235548.4]
  wire [5:0] _T_129; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235549.4]
  wire [5:0] _T_130; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235550.4]
  wire [5:0] _T_131; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235551.4]
  wire [5:0] _T_132; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235552.4]
  wire [5:0] _T_133; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235553.4]
  wire [126:0] _GEN_0; // @[rawFloatFromIN.scala 55:22:chipyard.TestHarness.RocketConfig.fir@235554.4]
  wire [126:0] _T_134; // @[rawFloatFromIN.scala 55:22:chipyard.TestHarness.RocketConfig.fir@235554.4]
  wire [5:0] _T_139; // @[rawFloatFromIN.scala 63:39:chipyard.TestHarness.RocketConfig.fir@235565.4]
  wire [7:0] _T_140; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@235566.4]
  RoundAnyRawFNToRecFN_1 roundAnyRawFNToRecFN ( // @[INToRecFN.scala 59:15:chipyard.TestHarness.RocketConfig.fir@235570.4]
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags)
  );
  assign intAsRawFloat_sign = io_signedIn & io_in[63]; // @[rawFloatFromIN.scala 50:29:chipyard.TestHarness.RocketConfig.fir@235421.4]
  assign _T_3 = 64'h0 - io_in; // @[rawFloatFromIN.scala 51:31:chipyard.TestHarness.RocketConfig.fir@235423.4]
  assign _T_4 = intAsRawFloat_sign ? _T_3 : io_in; // @[rawFloatFromIN.scala 51:24:chipyard.TestHarness.RocketConfig.fir@235424.4]
  assign _T_5 = {64'h0,_T_4}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@235425.4]
  assign _T_71 = _T_5[1] ? 6'h3e : 6'h3f; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235491.4]
  assign _T_72 = _T_5[2] ? 6'h3d : _T_71; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235492.4]
  assign _T_73 = _T_5[3] ? 6'h3c : _T_72; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235493.4]
  assign _T_74 = _T_5[4] ? 6'h3b : _T_73; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235494.4]
  assign _T_75 = _T_5[5] ? 6'h3a : _T_74; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235495.4]
  assign _T_76 = _T_5[6] ? 6'h39 : _T_75; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235496.4]
  assign _T_77 = _T_5[7] ? 6'h38 : _T_76; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235497.4]
  assign _T_78 = _T_5[8] ? 6'h37 : _T_77; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235498.4]
  assign _T_79 = _T_5[9] ? 6'h36 : _T_78; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235499.4]
  assign _T_80 = _T_5[10] ? 6'h35 : _T_79; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235500.4]
  assign _T_81 = _T_5[11] ? 6'h34 : _T_80; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235501.4]
  assign _T_82 = _T_5[12] ? 6'h33 : _T_81; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235502.4]
  assign _T_83 = _T_5[13] ? 6'h32 : _T_82; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235503.4]
  assign _T_84 = _T_5[14] ? 6'h31 : _T_83; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235504.4]
  assign _T_85 = _T_5[15] ? 6'h30 : _T_84; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235505.4]
  assign _T_86 = _T_5[16] ? 6'h2f : _T_85; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235506.4]
  assign _T_87 = _T_5[17] ? 6'h2e : _T_86; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235507.4]
  assign _T_88 = _T_5[18] ? 6'h2d : _T_87; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235508.4]
  assign _T_89 = _T_5[19] ? 6'h2c : _T_88; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235509.4]
  assign _T_90 = _T_5[20] ? 6'h2b : _T_89; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235510.4]
  assign _T_91 = _T_5[21] ? 6'h2a : _T_90; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235511.4]
  assign _T_92 = _T_5[22] ? 6'h29 : _T_91; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235512.4]
  assign _T_93 = _T_5[23] ? 6'h28 : _T_92; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235513.4]
  assign _T_94 = _T_5[24] ? 6'h27 : _T_93; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235514.4]
  assign _T_95 = _T_5[25] ? 6'h26 : _T_94; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235515.4]
  assign _T_96 = _T_5[26] ? 6'h25 : _T_95; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235516.4]
  assign _T_97 = _T_5[27] ? 6'h24 : _T_96; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235517.4]
  assign _T_98 = _T_5[28] ? 6'h23 : _T_97; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235518.4]
  assign _T_99 = _T_5[29] ? 6'h22 : _T_98; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235519.4]
  assign _T_100 = _T_5[30] ? 6'h21 : _T_99; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235520.4]
  assign _T_101 = _T_5[31] ? 6'h20 : _T_100; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235521.4]
  assign _T_102 = _T_5[32] ? 6'h1f : _T_101; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235522.4]
  assign _T_103 = _T_5[33] ? 6'h1e : _T_102; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235523.4]
  assign _T_104 = _T_5[34] ? 6'h1d : _T_103; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235524.4]
  assign _T_105 = _T_5[35] ? 6'h1c : _T_104; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235525.4]
  assign _T_106 = _T_5[36] ? 6'h1b : _T_105; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235526.4]
  assign _T_107 = _T_5[37] ? 6'h1a : _T_106; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235527.4]
  assign _T_108 = _T_5[38] ? 6'h19 : _T_107; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235528.4]
  assign _T_109 = _T_5[39] ? 6'h18 : _T_108; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235529.4]
  assign _T_110 = _T_5[40] ? 6'h17 : _T_109; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235530.4]
  assign _T_111 = _T_5[41] ? 6'h16 : _T_110; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235531.4]
  assign _T_112 = _T_5[42] ? 6'h15 : _T_111; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235532.4]
  assign _T_113 = _T_5[43] ? 6'h14 : _T_112; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235533.4]
  assign _T_114 = _T_5[44] ? 6'h13 : _T_113; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235534.4]
  assign _T_115 = _T_5[45] ? 6'h12 : _T_114; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235535.4]
  assign _T_116 = _T_5[46] ? 6'h11 : _T_115; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235536.4]
  assign _T_117 = _T_5[47] ? 6'h10 : _T_116; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235537.4]
  assign _T_118 = _T_5[48] ? 6'hf : _T_117; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235538.4]
  assign _T_119 = _T_5[49] ? 6'he : _T_118; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235539.4]
  assign _T_120 = _T_5[50] ? 6'hd : _T_119; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235540.4]
  assign _T_121 = _T_5[51] ? 6'hc : _T_120; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235541.4]
  assign _T_122 = _T_5[52] ? 6'hb : _T_121; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235542.4]
  assign _T_123 = _T_5[53] ? 6'ha : _T_122; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235543.4]
  assign _T_124 = _T_5[54] ? 6'h9 : _T_123; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235544.4]
  assign _T_125 = _T_5[55] ? 6'h8 : _T_124; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235545.4]
  assign _T_126 = _T_5[56] ? 6'h7 : _T_125; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235546.4]
  assign _T_127 = _T_5[57] ? 6'h6 : _T_126; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235547.4]
  assign _T_128 = _T_5[58] ? 6'h5 : _T_127; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235548.4]
  assign _T_129 = _T_5[59] ? 6'h4 : _T_128; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235549.4]
  assign _T_130 = _T_5[60] ? 6'h3 : _T_129; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235550.4]
  assign _T_131 = _T_5[61] ? 6'h2 : _T_130; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235551.4]
  assign _T_132 = _T_5[62] ? 6'h1 : _T_131; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235552.4]
  assign _T_133 = _T_5[63] ? 6'h0 : _T_132; // @[Mux.scala 47:69:chipyard.TestHarness.RocketConfig.fir@235553.4]
  assign _GEN_0 = {{63'd0}, _T_5[63:0]}; // @[rawFloatFromIN.scala 55:22:chipyard.TestHarness.RocketConfig.fir@235554.4]
  assign _T_134 = _GEN_0 << _T_133; // @[rawFloatFromIN.scala 55:22:chipyard.TestHarness.RocketConfig.fir@235554.4]
  assign _T_139 = ~_T_133; // @[rawFloatFromIN.scala 63:39:chipyard.TestHarness.RocketConfig.fir@235565.4]
  assign _T_140 = {2'h2,_T_139}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@235566.4]
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 72:23:chipyard.TestHarness.RocketConfig.fir@235577.4]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 73:23:chipyard.TestHarness.RocketConfig.fir@235578.4]
  assign roundAnyRawFNToRecFN_io_in_isZero = ~_T_134[63]; // @[INToRecFN.scala 69:44:chipyard.TestHarness.RocketConfig.fir@235574.4]
  assign roundAnyRawFNToRecFN_io_in_sign = io_signedIn & io_in[63]; // @[INToRecFN.scala 69:44:chipyard.TestHarness.RocketConfig.fir@235574.4]
  assign roundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(_T_140)}; // @[INToRecFN.scala 69:44:chipyard.TestHarness.RocketConfig.fir@235574.4]
  assign roundAnyRawFNToRecFN_io_in_sig = {{1'd0}, _T_134[63:0]}; // @[INToRecFN.scala 69:44:chipyard.TestHarness.RocketConfig.fir@235574.4]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[INToRecFN.scala 70:44:chipyard.TestHarness.RocketConfig.fir@235575.4]
endmodule
