module package_Anon( // @[:chipyard.TestHarness.RocketConfig.fir@195813.2]
  input  [19:0] io_x_ppn, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  input         io_x_u, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  input         io_x_ae, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  input         io_x_sw, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  input         io_x_sx, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  input         io_x_sr, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  input         io_x_pw, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  input         io_x_px, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  input         io_x_pr, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  input         io_x_pal, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  input         io_x_paa, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  input         io_x_eff, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  input         io_x_c, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  output [19:0] io_y_ppn, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  output        io_y_u, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  output        io_y_ae, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  output        io_y_sw, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  output        io_y_sx, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  output        io_y_sr, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  output        io_y_pw, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  output        io_y_px, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  output        io_y_pr, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  output        io_y_pal, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  output        io_y_paa, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  output        io_y_eff, // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
  output        io_y_c // @[:chipyard.TestHarness.RocketConfig.fir@195816.4]
);
  assign io_y_ppn = io_x_ppn; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@195821.4]
  assign io_y_u = io_x_u; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@195821.4]
  assign io_y_ae = io_x_ae; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@195821.4]
  assign io_y_sw = io_x_sw; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@195821.4]
  assign io_y_sx = io_x_sx; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@195821.4]
  assign io_y_sr = io_x_sr; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@195821.4]
  assign io_y_pw = io_x_pw; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@195821.4]
  assign io_y_px = io_x_px; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@195821.4]
  assign io_y_pr = io_x_pr; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@195821.4]
  assign io_y_pal = io_x_pal; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@195821.4]
  assign io_y_paa = io_x_paa; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@195821.4]
  assign io_y_eff = io_x_eff; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@195821.4]
  assign io_y_c = io_x_c; // @[package.scala 218:12:chipyard.TestHarness.RocketConfig.fir@195821.4]
endmodule
