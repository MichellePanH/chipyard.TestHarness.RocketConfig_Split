module DCacheModuleImpl_Anon_1( // @[:chipyard.TestHarness.RocketConfig.fir@213366.2]
  input         io_in_0_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [39:0] io_in_0_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [5:0]  io_in_0_bits_idx, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [21:0] io_in_0_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input         io_in_1_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [39:0] io_in_1_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [5:0]  io_in_1_bits_idx, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [21:0] io_in_1_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input         io_in_2_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [39:0] io_in_2_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [5:0]  io_in_2_bits_idx, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [3:0]  io_in_2_bits_way_en, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [21:0] io_in_2_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input         io_in_3_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [39:0] io_in_3_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [5:0]  io_in_3_bits_idx, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [3:0]  io_in_3_bits_way_en, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [21:0] io_in_3_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  output        io_in_4_ready, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input         io_in_4_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [39:0] io_in_4_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [5:0]  io_in_4_bits_idx, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [3:0]  io_in_4_bits_way_en, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [21:0] io_in_4_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  output        io_in_5_ready, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input         io_in_5_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [39:0] io_in_5_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [5:0]  io_in_5_bits_idx, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  output        io_in_6_ready, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input         io_in_6_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [39:0] io_in_6_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [5:0]  io_in_6_bits_idx, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [3:0]  io_in_6_bits_way_en, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [21:0] io_in_6_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  output        io_in_7_ready, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input         io_in_7_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [39:0] io_in_7_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [5:0]  io_in_7_bits_idx, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [3:0]  io_in_7_bits_way_en, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  input  [21:0] io_in_7_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  output        io_out_valid, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  output        io_out_bits_write, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  output [39:0] io_out_bits_addr, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  output [5:0]  io_out_bits_idx, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  output [3:0]  io_out_bits_way_en, // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
  output [21:0] io_out_bits_data // @[:chipyard.TestHarness.RocketConfig.fir@213369.4]
);
  wire [21:0] _GEN_1; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213377.4]
  wire [3:0] _GEN_2; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213377.4]
  wire [5:0] _GEN_3; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213377.4]
  wire [39:0] _GEN_4; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213377.4]
  wire [21:0] _GEN_13; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213393.4]
  wire [3:0] _GEN_14; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213393.4]
  wire [5:0] _GEN_15; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213393.4]
  wire [39:0] _GEN_16; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213393.4]
  wire [21:0] _GEN_19; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213401.4]
  wire [3:0] _GEN_20; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213401.4]
  wire [5:0] _GEN_21; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213401.4]
  wire [39:0] _GEN_22; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213401.4]
  wire  _GEN_23; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213401.4]
  wire [21:0] _GEN_25; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213409.4]
  wire [3:0] _GEN_26; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213409.4]
  wire [5:0] _GEN_27; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213409.4]
  wire [39:0] _GEN_28; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213409.4]
  wire  _GEN_29; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213409.4]
  wire [21:0] _GEN_31; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213417.4]
  wire [3:0] _GEN_32; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213417.4]
  wire [5:0] _GEN_33; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213417.4]
  wire [39:0] _GEN_34; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213417.4]
  wire  _GEN_35; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213417.4]
  wire  _T; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213433.4]
  wire  _T_1; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213434.4]
  wire  _T_2; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213435.4]
  wire  _T_3; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213436.4]
  wire  _T_5; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213438.4]
  wire  grant_7; // @[Arbiter.scala 31:78:chipyard.TestHarness.RocketConfig.fir@213445.4]
  wire  _T_14; // @[Arbiter.scala 135:19:chipyard.TestHarness.RocketConfig.fir@213462.4]
  assign _GEN_1 = io_in_6_valid ? io_in_6_bits_data : io_in_7_bits_data; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213377.4]
  assign _GEN_2 = io_in_6_valid ? io_in_6_bits_way_en : io_in_7_bits_way_en; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213377.4]
  assign _GEN_3 = io_in_6_valid ? io_in_6_bits_idx : io_in_7_bits_idx; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213377.4]
  assign _GEN_4 = io_in_6_valid ? io_in_6_bits_addr : io_in_7_bits_addr; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213377.4]
  assign _GEN_13 = io_in_4_valid ? io_in_4_bits_data : _GEN_1; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213393.4]
  assign _GEN_14 = io_in_4_valid ? io_in_4_bits_way_en : _GEN_2; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213393.4]
  assign _GEN_15 = io_in_4_valid ? io_in_4_bits_idx : _GEN_3; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213393.4]
  assign _GEN_16 = io_in_4_valid ? io_in_4_bits_addr : _GEN_4; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213393.4]
  assign _GEN_19 = io_in_3_valid ? io_in_3_bits_data : _GEN_13; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213401.4]
  assign _GEN_20 = io_in_3_valid ? io_in_3_bits_way_en : _GEN_14; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213401.4]
  assign _GEN_21 = io_in_3_valid ? io_in_3_bits_idx : _GEN_15; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213401.4]
  assign _GEN_22 = io_in_3_valid ? io_in_3_bits_addr : _GEN_16; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213401.4]
  assign _GEN_23 = io_in_3_valid | io_in_4_valid; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213401.4]
  assign _GEN_25 = io_in_2_valid ? io_in_2_bits_data : _GEN_19; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213409.4]
  assign _GEN_26 = io_in_2_valid ? io_in_2_bits_way_en : _GEN_20; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213409.4]
  assign _GEN_27 = io_in_2_valid ? io_in_2_bits_idx : _GEN_21; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213409.4]
  assign _GEN_28 = io_in_2_valid ? io_in_2_bits_addr : _GEN_22; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213409.4]
  assign _GEN_29 = io_in_2_valid | _GEN_23; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213409.4]
  assign _GEN_31 = io_in_1_valid ? io_in_1_bits_data : _GEN_25; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213417.4]
  assign _GEN_32 = io_in_1_valid ? 4'h0 : _GEN_26; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213417.4]
  assign _GEN_33 = io_in_1_valid ? io_in_1_bits_idx : _GEN_27; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213417.4]
  assign _GEN_34 = io_in_1_valid ? io_in_1_bits_addr : _GEN_28; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213417.4]
  assign _GEN_35 = io_in_1_valid | _GEN_29; // @[Arbiter.scala 126:27:chipyard.TestHarness.RocketConfig.fir@213417.4]
  assign _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213433.4]
  assign _T_1 = _T | io_in_2_valid; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213434.4]
  assign _T_2 = _T_1 | io_in_3_valid; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213435.4]
  assign _T_3 = _T_2 | io_in_4_valid; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213436.4]
  assign _T_5 = _T_3 | io_in_6_valid; // @[Arbiter.scala 31:68:chipyard.TestHarness.RocketConfig.fir@213438.4]
  assign grant_7 = ~_T_5; // @[Arbiter.scala 31:78:chipyard.TestHarness.RocketConfig.fir@213445.4]
  assign _T_14 = ~grant_7; // @[Arbiter.scala 135:19:chipyard.TestHarness.RocketConfig.fir@213462.4]
  assign io_in_4_ready = ~_T_2; // @[Arbiter.scala 134:14:chipyard.TestHarness.RocketConfig.fir@213455.4]
  assign io_in_5_ready = ~_T_3; // @[Arbiter.scala 134:14:chipyard.TestHarness.RocketConfig.fir@213457.4]
  assign io_in_6_ready = ~_T_3; // @[Arbiter.scala 134:14:chipyard.TestHarness.RocketConfig.fir@213459.4]
  assign io_in_7_ready = ~_T_5; // @[Arbiter.scala 134:14:chipyard.TestHarness.RocketConfig.fir@213461.4]
  assign io_out_valid = _T_14 | io_in_7_valid; // @[Arbiter.scala 135:16:chipyard.TestHarness.RocketConfig.fir@213464.4]
  assign io_out_bits_write = io_in_0_valid | _GEN_35; // @[Arbiter.scala 124:15:chipyard.TestHarness.RocketConfig.fir@213376.4 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213383.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213391.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213399.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213407.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213415.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213423.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213431.6]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_34; // @[Arbiter.scala 124:15:chipyard.TestHarness.RocketConfig.fir@213375.4 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213382.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213390.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213398.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213406.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213414.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213422.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213430.6]
  assign io_out_bits_idx = io_in_0_valid ? io_in_0_bits_idx : _GEN_33; // @[Arbiter.scala 124:15:chipyard.TestHarness.RocketConfig.fir@213374.4 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213381.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213389.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213397.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213405.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213413.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213421.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213429.6]
  assign io_out_bits_way_en = io_in_0_valid ? 4'hf : _GEN_32; // @[Arbiter.scala 124:15:chipyard.TestHarness.RocketConfig.fir@213373.4 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213380.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213388.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213396.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213404.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213412.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213420.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213428.6]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : _GEN_31; // @[Arbiter.scala 124:15:chipyard.TestHarness.RocketConfig.fir@213372.4 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213379.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213387.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213395.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213403.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213411.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213419.6 Arbiter.scala 128:19:chipyard.TestHarness.RocketConfig.fir@213427.6]
endmodule
