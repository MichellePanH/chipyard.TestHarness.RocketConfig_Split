module Scheduler( // @[:chipyard.TestHarness.RocketConfig.fir@100021.2]
  input         clock, // @[:chipyard.TestHarness.RocketConfig.fir@100022.4]
  input         reset, // @[:chipyard.TestHarness.RocketConfig.fir@100023.4]
  output        io_in_a_ready, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_in_a_valid, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [2:0]  io_in_a_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [2:0]  io_in_a_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [2:0]  io_in_a_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [2:0]  io_in_a_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [31:0] io_in_a_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [7:0]  io_in_a_bits_mask, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [63:0] io_in_a_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_in_a_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_in_b_ready, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output        io_in_b_valid, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [1:0]  io_in_b_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [31:0] io_in_b_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output        io_in_c_ready, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_in_c_valid, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [2:0]  io_in_c_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [2:0]  io_in_c_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [2:0]  io_in_c_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [2:0]  io_in_c_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [31:0] io_in_c_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [63:0] io_in_c_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_in_c_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_in_d_ready, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output        io_in_d_valid, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [2:0]  io_in_d_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [1:0]  io_in_d_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [2:0]  io_in_d_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [2:0]  io_in_d_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [2:0]  io_in_d_bits_sink, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output        io_in_d_bits_denied, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [63:0] io_in_d_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output        io_in_d_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_in_e_valid, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [2:0]  io_in_e_bits_sink, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_out_a_ready, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output        io_out_a_valid, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [2:0]  io_out_a_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [2:0]  io_out_a_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [2:0]  io_out_a_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [2:0]  io_out_a_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [31:0] io_out_a_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [7:0]  io_out_a_bits_mask, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [63:0] io_out_a_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output        io_out_a_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_out_c_ready, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output        io_out_c_valid, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [2:0]  io_out_c_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [2:0]  io_out_c_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [2:0]  io_out_c_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [2:0]  io_out_c_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [31:0] io_out_c_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [63:0] io_out_c_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output        io_out_c_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output        io_out_d_ready, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_out_d_valid, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [2:0]  io_out_d_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [1:0]  io_out_d_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [2:0]  io_out_d_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [2:0]  io_out_d_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [2:0]  io_out_d_bits_sink, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_out_d_bits_denied, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [63:0] io_out_d_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_out_d_bits_corrupt, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output        io_out_e_valid, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output [2:0]  io_out_e_bits_sink, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output        io_req_ready, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_req_valid, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input  [31:0] io_req_bits_address, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  input         io_resp_ready, // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
  output        io_resp_valid // @[:chipyard.TestHarness.RocketConfig.fir@100024.4]
);
  wire  sourceA_clock; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire  sourceA_reset; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire  sourceA_io_req_ready; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire  sourceA_io_req_valid; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire [11:0] sourceA_io_req_bits_tag; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire [9:0] sourceA_io_req_bits_set; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire [2:0] sourceA_io_req_bits_param; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire [2:0] sourceA_io_req_bits_source; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire  sourceA_io_req_bits_block; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire  sourceA_io_a_ready; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire  sourceA_io_a_valid; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire [2:0] sourceA_io_a_bits_opcode; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire [2:0] sourceA_io_a_bits_param; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire [2:0] sourceA_io_a_bits_size; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire [2:0] sourceA_io_a_bits_source; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire [31:0] sourceA_io_a_bits_address; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire [7:0] sourceA_io_a_bits_mask; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire [63:0] sourceA_io_a_bits_data; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire  sourceA_io_a_bits_corrupt; // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
  wire  sourceB_clock; // @[Scheduler.scala 39:23:chipyard.TestHarness.RocketConfig.fir@100033.4]
  wire  sourceB_reset; // @[Scheduler.scala 39:23:chipyard.TestHarness.RocketConfig.fir@100033.4]
  wire  sourceB_io_req_ready; // @[Scheduler.scala 39:23:chipyard.TestHarness.RocketConfig.fir@100033.4]
  wire  sourceB_io_req_valid; // @[Scheduler.scala 39:23:chipyard.TestHarness.RocketConfig.fir@100033.4]
  wire [2:0] sourceB_io_req_bits_param; // @[Scheduler.scala 39:23:chipyard.TestHarness.RocketConfig.fir@100033.4]
  wire [11:0] sourceB_io_req_bits_tag; // @[Scheduler.scala 39:23:chipyard.TestHarness.RocketConfig.fir@100033.4]
  wire [9:0] sourceB_io_req_bits_set; // @[Scheduler.scala 39:23:chipyard.TestHarness.RocketConfig.fir@100033.4]
  wire  sourceB_io_req_bits_clients; // @[Scheduler.scala 39:23:chipyard.TestHarness.RocketConfig.fir@100033.4]
  wire  sourceB_io_b_ready; // @[Scheduler.scala 39:23:chipyard.TestHarness.RocketConfig.fir@100033.4]
  wire  sourceB_io_b_valid; // @[Scheduler.scala 39:23:chipyard.TestHarness.RocketConfig.fir@100033.4]
  wire [1:0] sourceB_io_b_bits_param; // @[Scheduler.scala 39:23:chipyard.TestHarness.RocketConfig.fir@100033.4]
  wire [31:0] sourceB_io_b_bits_address; // @[Scheduler.scala 39:23:chipyard.TestHarness.RocketConfig.fir@100033.4]
  wire  sourceC_clock; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire  sourceC_reset; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire  sourceC_io_req_ready; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire  sourceC_io_req_valid; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [2:0] sourceC_io_req_bits_opcode; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [2:0] sourceC_io_req_bits_param; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [2:0] sourceC_io_req_bits_source; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [11:0] sourceC_io_req_bits_tag; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [9:0] sourceC_io_req_bits_set; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [2:0] sourceC_io_req_bits_way; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire  sourceC_io_req_bits_dirty; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire  sourceC_io_c_ready; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire  sourceC_io_c_valid; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [2:0] sourceC_io_c_bits_opcode; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [2:0] sourceC_io_c_bits_param; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [2:0] sourceC_io_c_bits_size; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [2:0] sourceC_io_c_bits_source; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [31:0] sourceC_io_c_bits_address; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [63:0] sourceC_io_c_bits_data; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire  sourceC_io_c_bits_corrupt; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire  sourceC_io_bs_adr_ready; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire  sourceC_io_bs_adr_valid; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [2:0] sourceC_io_bs_adr_bits_way; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [9:0] sourceC_io_bs_adr_bits_set; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [2:0] sourceC_io_bs_adr_bits_beat; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [63:0] sourceC_io_bs_dat_data; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [9:0] sourceC_io_evict_req_set; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire [2:0] sourceC_io_evict_req_way; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire  sourceC_io_evict_safe; // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
  wire  sourceD_clock; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_reset; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_req_ready; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_req_valid; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_req_bits_prio_0; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_req_bits_prio_2; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_req_bits_opcode; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_req_bits_param; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_req_bits_size; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_req_bits_source; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [5:0] sourceD_io_req_bits_offset; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [5:0] sourceD_io_req_bits_put; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [9:0] sourceD_io_req_bits_set; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_req_bits_sink; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_req_bits_way; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_req_bits_bad; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_d_ready; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_d_valid; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_d_bits_opcode; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [1:0] sourceD_io_d_bits_param; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_d_bits_size; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_d_bits_source; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_d_bits_sink; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_d_bits_denied; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [63:0] sourceD_io_d_bits_data; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_d_bits_corrupt; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_pb_pop_ready; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_pb_pop_valid; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [5:0] sourceD_io_pb_pop_bits_index; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_pb_pop_bits_last; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [63:0] sourceD_io_pb_beat_data; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [7:0] sourceD_io_pb_beat_mask; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_pb_beat_corrupt; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_rel_pop_ready; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_rel_pop_valid; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [5:0] sourceD_io_rel_pop_bits_index; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_rel_pop_bits_last; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [63:0] sourceD_io_rel_beat_data; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_rel_beat_corrupt; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_bs_radr_ready; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_bs_radr_valid; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_bs_radr_bits_way; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [9:0] sourceD_io_bs_radr_bits_set; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_bs_radr_bits_beat; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_bs_radr_bits_mask; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [63:0] sourceD_io_bs_rdat_data; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_bs_wadr_ready; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_bs_wadr_valid; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_bs_wadr_bits_way; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [9:0] sourceD_io_bs_wadr_bits_set; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_bs_wadr_bits_beat; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_bs_wadr_bits_mask; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [63:0] sourceD_io_bs_wdat_data; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [9:0] sourceD_io_evict_req_set; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_evict_req_way; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_evict_safe; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [9:0] sourceD_io_grant_req_set; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire [2:0] sourceD_io_grant_req_way; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceD_io_grant_safe; // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
  wire  sourceE_clock; // @[Scheduler.scala 42:23:chipyard.TestHarness.RocketConfig.fir@100045.4]
  wire  sourceE_reset; // @[Scheduler.scala 42:23:chipyard.TestHarness.RocketConfig.fir@100045.4]
  wire  sourceE_io_req_ready; // @[Scheduler.scala 42:23:chipyard.TestHarness.RocketConfig.fir@100045.4]
  wire  sourceE_io_req_valid; // @[Scheduler.scala 42:23:chipyard.TestHarness.RocketConfig.fir@100045.4]
  wire [2:0] sourceE_io_req_bits_sink; // @[Scheduler.scala 42:23:chipyard.TestHarness.RocketConfig.fir@100045.4]
  wire  sourceE_io_e_valid; // @[Scheduler.scala 42:23:chipyard.TestHarness.RocketConfig.fir@100045.4]
  wire [2:0] sourceE_io_e_bits_sink; // @[Scheduler.scala 42:23:chipyard.TestHarness.RocketConfig.fir@100045.4]
  wire  sourceX_clock; // @[Scheduler.scala 43:23:chipyard.TestHarness.RocketConfig.fir@100049.4]
  wire  sourceX_reset; // @[Scheduler.scala 43:23:chipyard.TestHarness.RocketConfig.fir@100049.4]
  wire  sourceX_io_req_ready; // @[Scheduler.scala 43:23:chipyard.TestHarness.RocketConfig.fir@100049.4]
  wire  sourceX_io_req_valid; // @[Scheduler.scala 43:23:chipyard.TestHarness.RocketConfig.fir@100049.4]
  wire  sourceX_io_x_ready; // @[Scheduler.scala 43:23:chipyard.TestHarness.RocketConfig.fir@100049.4]
  wire  sourceX_io_x_valid; // @[Scheduler.scala 43:23:chipyard.TestHarness.RocketConfig.fir@100049.4]
  wire  sinkA_clock; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire  sinkA_reset; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire  sinkA_io_req_ready; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire  sinkA_io_req_valid; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [2:0] sinkA_io_req_bits_opcode; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [2:0] sinkA_io_req_bits_param; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [2:0] sinkA_io_req_bits_size; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [2:0] sinkA_io_req_bits_source; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [11:0] sinkA_io_req_bits_tag; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [5:0] sinkA_io_req_bits_offset; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [5:0] sinkA_io_req_bits_put; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [9:0] sinkA_io_req_bits_set; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire  sinkA_io_a_ready; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire  sinkA_io_a_valid; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [2:0] sinkA_io_a_bits_opcode; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [2:0] sinkA_io_a_bits_param; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [2:0] sinkA_io_a_bits_size; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [2:0] sinkA_io_a_bits_source; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [31:0] sinkA_io_a_bits_address; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [7:0] sinkA_io_a_bits_mask; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [63:0] sinkA_io_a_bits_data; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire  sinkA_io_a_bits_corrupt; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire  sinkA_io_pb_pop_ready; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire  sinkA_io_pb_pop_valid; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [5:0] sinkA_io_pb_pop_bits_index; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire  sinkA_io_pb_pop_bits_last; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [63:0] sinkA_io_pb_beat_data; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire [7:0] sinkA_io_pb_beat_mask; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire  sinkA_io_pb_beat_corrupt; // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
  wire  sinkC_clock; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_reset; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_req_ready; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_req_valid; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [2:0] sinkC_io_req_bits_opcode; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [2:0] sinkC_io_req_bits_param; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [2:0] sinkC_io_req_bits_size; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [2:0] sinkC_io_req_bits_source; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [11:0] sinkC_io_req_bits_tag; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [5:0] sinkC_io_req_bits_offset; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [5:0] sinkC_io_req_bits_put; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [9:0] sinkC_io_req_bits_set; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_resp_valid; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_resp_bits_last; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [9:0] sinkC_io_resp_bits_set; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [11:0] sinkC_io_resp_bits_tag; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [2:0] sinkC_io_resp_bits_source; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [2:0] sinkC_io_resp_bits_param; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_resp_bits_data; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_c_ready; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_c_valid; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [2:0] sinkC_io_c_bits_opcode; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [2:0] sinkC_io_c_bits_param; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [2:0] sinkC_io_c_bits_size; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [2:0] sinkC_io_c_bits_source; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [31:0] sinkC_io_c_bits_address; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [63:0] sinkC_io_c_bits_data; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_c_bits_corrupt; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [9:0] sinkC_io_set; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [2:0] sinkC_io_way; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_bs_adr_ready; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_bs_adr_valid; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_bs_adr_bits_noop; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [2:0] sinkC_io_bs_adr_bits_way; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [9:0] sinkC_io_bs_adr_bits_set; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [2:0] sinkC_io_bs_adr_bits_beat; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_bs_adr_bits_mask; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [63:0] sinkC_io_bs_dat_data; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_rel_pop_ready; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_rel_pop_valid; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [5:0] sinkC_io_rel_pop_bits_index; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_rel_pop_bits_last; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire [63:0] sinkC_io_rel_beat_data; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkC_io_rel_beat_corrupt; // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
  wire  sinkD_clock; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire  sinkD_reset; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire  sinkD_io_resp_valid; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire  sinkD_io_resp_bits_last; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [2:0] sinkD_io_resp_bits_opcode; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [2:0] sinkD_io_resp_bits_param; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [2:0] sinkD_io_resp_bits_source; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [2:0] sinkD_io_resp_bits_sink; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire  sinkD_io_resp_bits_denied; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire  sinkD_io_d_ready; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire  sinkD_io_d_valid; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [2:0] sinkD_io_d_bits_opcode; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [1:0] sinkD_io_d_bits_param; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [2:0] sinkD_io_d_bits_size; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [2:0] sinkD_io_d_bits_source; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [2:0] sinkD_io_d_bits_sink; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire  sinkD_io_d_bits_denied; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [63:0] sinkD_io_d_bits_data; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire  sinkD_io_d_bits_corrupt; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [2:0] sinkD_io_source; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [2:0] sinkD_io_way; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [9:0] sinkD_io_set; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire  sinkD_io_bs_adr_ready; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire  sinkD_io_bs_adr_valid; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire  sinkD_io_bs_adr_bits_noop; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [2:0] sinkD_io_bs_adr_bits_way; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [9:0] sinkD_io_bs_adr_bits_set; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [2:0] sinkD_io_bs_adr_bits_beat; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [63:0] sinkD_io_bs_dat_data; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [9:0] sinkD_io_grant_req_set; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire [2:0] sinkD_io_grant_req_way; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire  sinkD_io_grant_safe; // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
  wire  sinkE_io_resp_valid; // @[Scheduler.scala 55:21:chipyard.TestHarness.RocketConfig.fir@100071.4]
  wire [2:0] sinkE_io_resp_bits_sink; // @[Scheduler.scala 55:21:chipyard.TestHarness.RocketConfig.fir@100071.4]
  wire  sinkE_io_e_valid; // @[Scheduler.scala 55:21:chipyard.TestHarness.RocketConfig.fir@100071.4]
  wire [2:0] sinkE_io_e_bits_sink; // @[Scheduler.scala 55:21:chipyard.TestHarness.RocketConfig.fir@100071.4]
  wire  sinkX_clock; // @[Scheduler.scala 56:21:chipyard.TestHarness.RocketConfig.fir@100075.4]
  wire  sinkX_reset; // @[Scheduler.scala 56:21:chipyard.TestHarness.RocketConfig.fir@100075.4]
  wire  sinkX_io_req_ready; // @[Scheduler.scala 56:21:chipyard.TestHarness.RocketConfig.fir@100075.4]
  wire  sinkX_io_req_valid; // @[Scheduler.scala 56:21:chipyard.TestHarness.RocketConfig.fir@100075.4]
  wire [11:0] sinkX_io_req_bits_tag; // @[Scheduler.scala 56:21:chipyard.TestHarness.RocketConfig.fir@100075.4]
  wire [9:0] sinkX_io_req_bits_set; // @[Scheduler.scala 56:21:chipyard.TestHarness.RocketConfig.fir@100075.4]
  wire  sinkX_io_x_ready; // @[Scheduler.scala 56:21:chipyard.TestHarness.RocketConfig.fir@100075.4]
  wire  sinkX_io_x_valid; // @[Scheduler.scala 56:21:chipyard.TestHarness.RocketConfig.fir@100075.4]
  wire [31:0] sinkX_io_x_bits_address; // @[Scheduler.scala 56:21:chipyard.TestHarness.RocketConfig.fir@100075.4]
  wire  directory_clock; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire  directory_reset; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire  directory_io_write_ready; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire  directory_io_write_valid; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire [9:0] directory_io_write_bits_set; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire [2:0] directory_io_write_bits_way; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire  directory_io_write_bits_data_dirty; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire [1:0] directory_io_write_bits_data_state; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire  directory_io_write_bits_data_clients; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire [11:0] directory_io_write_bits_data_tag; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire  directory_io_read_valid; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire [9:0] directory_io_read_bits_set; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire [11:0] directory_io_read_bits_tag; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire  directory_io_result_bits_dirty; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire [1:0] directory_io_result_bits_state; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire  directory_io_result_bits_clients; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire [11:0] directory_io_result_bits_tag; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire  directory_io_result_bits_hit; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire [2:0] directory_io_result_bits_way; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire  directory_io_ready; // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
  wire  bankedStore_clock; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sinkC_adr_ready; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sinkC_adr_valid; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sinkC_adr_bits_noop; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [2:0] bankedStore_io_sinkC_adr_bits_way; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [9:0] bankedStore_io_sinkC_adr_bits_set; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [2:0] bankedStore_io_sinkC_adr_bits_beat; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sinkC_adr_bits_mask; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [63:0] bankedStore_io_sinkC_dat_data; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sinkD_adr_ready; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sinkD_adr_valid; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sinkD_adr_bits_noop; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [2:0] bankedStore_io_sinkD_adr_bits_way; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [9:0] bankedStore_io_sinkD_adr_bits_set; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [2:0] bankedStore_io_sinkD_adr_bits_beat; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [63:0] bankedStore_io_sinkD_dat_data; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sourceC_adr_ready; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sourceC_adr_valid; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [2:0] bankedStore_io_sourceC_adr_bits_way; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [9:0] bankedStore_io_sourceC_adr_bits_set; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [2:0] bankedStore_io_sourceC_adr_bits_beat; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [63:0] bankedStore_io_sourceC_dat_data; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sourceD_radr_ready; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sourceD_radr_valid; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [2:0] bankedStore_io_sourceD_radr_bits_way; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [9:0] bankedStore_io_sourceD_radr_bits_set; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [2:0] bankedStore_io_sourceD_radr_bits_beat; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sourceD_radr_bits_mask; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [63:0] bankedStore_io_sourceD_rdat_data; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sourceD_wadr_ready; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sourceD_wadr_valid; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [2:0] bankedStore_io_sourceD_wadr_bits_way; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [9:0] bankedStore_io_sourceD_wadr_bits_set; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [2:0] bankedStore_io_sourceD_wadr_bits_beat; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  bankedStore_io_sourceD_wadr_bits_mask; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire [63:0] bankedStore_io_sourceD_wdat_data; // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
  wire  requests_clock; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire  requests_reset; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire  requests_io_push_ready; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire  requests_io_push_valid; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [4:0] requests_io_push_bits_index; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire  requests_io_push_bits_data_prio_0; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire  requests_io_push_bits_data_prio_2; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire  requests_io_push_bits_data_control; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [2:0] requests_io_push_bits_data_opcode; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [2:0] requests_io_push_bits_data_param; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [2:0] requests_io_push_bits_data_size; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [2:0] requests_io_push_bits_data_source; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [11:0] requests_io_push_bits_data_tag; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [5:0] requests_io_push_bits_data_offset; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [5:0] requests_io_push_bits_data_put; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [20:0] requests_io_valid; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire  requests_io_pop_valid; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [4:0] requests_io_pop_bits; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire  requests_io_data_prio_0; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire  requests_io_data_prio_1; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire  requests_io_data_prio_2; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire  requests_io_data_control; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [2:0] requests_io_data_opcode; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [2:0] requests_io_data_param; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [2:0] requests_io_data_size; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [2:0] requests_io_data_source; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [11:0] requests_io_data_tag; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [5:0] requests_io_data_offset; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire [5:0] requests_io_data_put; // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
  wire  abc_mshrs_0_clock; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_reset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_allocate_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_allocate_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_allocate_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_allocate_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_allocate_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_allocate_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_allocate_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_allocate_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_allocate_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [11:0] abc_mshrs_0_io_allocate_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [5:0] abc_mshrs_0_io_allocate_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [5:0] abc_mshrs_0_io_allocate_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [9:0] abc_mshrs_0_io_allocate_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_allocate_bits_repeat; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_directory_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_directory_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [1:0] abc_mshrs_0_io_directory_bits_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_directory_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [11:0] abc_mshrs_0_io_directory_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_directory_bits_hit; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_directory_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_status_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [9:0] abc_mshrs_0_io_status_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [11:0] abc_mshrs_0_io_status_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_status_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_status_bits_blockB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_status_bits_nestB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_status_bits_blockC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_status_bits_nestC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_ready; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_a_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [11:0] abc_mshrs_0_io_schedule_bits_a_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [9:0] abc_mshrs_0_io_schedule_bits_a_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_schedule_bits_a_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_a_bits_block; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_b_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_schedule_bits_b_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [11:0] abc_mshrs_0_io_schedule_bits_b_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [9:0] abc_mshrs_0_io_schedule_bits_b_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_b_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_c_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_schedule_bits_c_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_schedule_bits_c_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [11:0] abc_mshrs_0_io_schedule_bits_c_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [9:0] abc_mshrs_0_io_schedule_bits_c_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_schedule_bits_c_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_c_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_d_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_d_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_d_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_d_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_d_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_schedule_bits_d_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_schedule_bits_d_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_schedule_bits_d_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_schedule_bits_d_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [11:0] abc_mshrs_0_io_schedule_bits_d_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [5:0] abc_mshrs_0_io_schedule_bits_d_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [5:0] abc_mshrs_0_io_schedule_bits_d_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [9:0] abc_mshrs_0_io_schedule_bits_d_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_schedule_bits_d_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_d_bits_bad; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_e_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_schedule_bits_e_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_x_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_dir_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [9:0] abc_mshrs_0_io_schedule_bits_dir_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_schedule_bits_dir_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [1:0] abc_mshrs_0_io_schedule_bits_dir_bits_data_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_dir_bits_data_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [11:0] abc_mshrs_0_io_schedule_bits_dir_bits_data_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_schedule_bits_reload; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_sinkc_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_sinkc_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [11:0] abc_mshrs_0_io_sinkc_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_sinkc_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_sinkc_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_sinkc_bits_data; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_sinkd_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_sinkd_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_sinkd_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_sinkd_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [2:0] abc_mshrs_0_io_sinkd_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_sinkd_bits_denied; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_sinke_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [9:0] abc_mshrs_0_io_nestedwb_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire [11:0] abc_mshrs_0_io_nestedwb_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_nestedwb_b_toN; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_nestedwb_b_toB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_nestedwb_b_clr_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_0_io_nestedwb_c_set_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
  wire  abc_mshrs_1_clock; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_reset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_allocate_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_allocate_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_allocate_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_allocate_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_allocate_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_allocate_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_allocate_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_allocate_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_allocate_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [11:0] abc_mshrs_1_io_allocate_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [5:0] abc_mshrs_1_io_allocate_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [5:0] abc_mshrs_1_io_allocate_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [9:0] abc_mshrs_1_io_allocate_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_allocate_bits_repeat; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_directory_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_directory_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [1:0] abc_mshrs_1_io_directory_bits_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_directory_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [11:0] abc_mshrs_1_io_directory_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_directory_bits_hit; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_directory_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_status_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [9:0] abc_mshrs_1_io_status_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [11:0] abc_mshrs_1_io_status_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_status_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_status_bits_blockB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_status_bits_nestB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_status_bits_blockC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_status_bits_nestC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_ready; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_a_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [11:0] abc_mshrs_1_io_schedule_bits_a_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [9:0] abc_mshrs_1_io_schedule_bits_a_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_schedule_bits_a_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_a_bits_block; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_b_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_schedule_bits_b_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [11:0] abc_mshrs_1_io_schedule_bits_b_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [9:0] abc_mshrs_1_io_schedule_bits_b_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_b_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_c_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_schedule_bits_c_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_schedule_bits_c_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [11:0] abc_mshrs_1_io_schedule_bits_c_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [9:0] abc_mshrs_1_io_schedule_bits_c_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_schedule_bits_c_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_c_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_d_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_d_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_d_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_d_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_d_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_schedule_bits_d_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_schedule_bits_d_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_schedule_bits_d_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_schedule_bits_d_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [11:0] abc_mshrs_1_io_schedule_bits_d_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [5:0] abc_mshrs_1_io_schedule_bits_d_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [5:0] abc_mshrs_1_io_schedule_bits_d_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [9:0] abc_mshrs_1_io_schedule_bits_d_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_schedule_bits_d_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_d_bits_bad; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_e_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_schedule_bits_e_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_x_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_dir_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [9:0] abc_mshrs_1_io_schedule_bits_dir_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_schedule_bits_dir_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [1:0] abc_mshrs_1_io_schedule_bits_dir_bits_data_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_dir_bits_data_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [11:0] abc_mshrs_1_io_schedule_bits_dir_bits_data_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_schedule_bits_reload; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_sinkc_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_sinkc_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [11:0] abc_mshrs_1_io_sinkc_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_sinkc_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_sinkc_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_sinkc_bits_data; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_sinkd_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_sinkd_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_sinkd_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_sinkd_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [2:0] abc_mshrs_1_io_sinkd_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_sinkd_bits_denied; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_sinke_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [9:0] abc_mshrs_1_io_nestedwb_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire [11:0] abc_mshrs_1_io_nestedwb_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_nestedwb_b_toN; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_nestedwb_b_toB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_nestedwb_b_clr_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_1_io_nestedwb_c_set_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
  wire  abc_mshrs_2_clock; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_reset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_allocate_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_allocate_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_allocate_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_allocate_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_allocate_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_allocate_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_allocate_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_allocate_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_allocate_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [11:0] abc_mshrs_2_io_allocate_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [5:0] abc_mshrs_2_io_allocate_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [5:0] abc_mshrs_2_io_allocate_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [9:0] abc_mshrs_2_io_allocate_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_allocate_bits_repeat; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_directory_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_directory_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [1:0] abc_mshrs_2_io_directory_bits_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_directory_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [11:0] abc_mshrs_2_io_directory_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_directory_bits_hit; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_directory_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_status_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [9:0] abc_mshrs_2_io_status_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [11:0] abc_mshrs_2_io_status_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_status_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_status_bits_blockB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_status_bits_nestB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_status_bits_blockC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_status_bits_nestC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_ready; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_a_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [11:0] abc_mshrs_2_io_schedule_bits_a_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [9:0] abc_mshrs_2_io_schedule_bits_a_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_schedule_bits_a_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_a_bits_block; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_b_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_schedule_bits_b_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [11:0] abc_mshrs_2_io_schedule_bits_b_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [9:0] abc_mshrs_2_io_schedule_bits_b_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_b_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_c_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_schedule_bits_c_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_schedule_bits_c_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [11:0] abc_mshrs_2_io_schedule_bits_c_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [9:0] abc_mshrs_2_io_schedule_bits_c_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_schedule_bits_c_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_c_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_d_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_d_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_d_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_d_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_d_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_schedule_bits_d_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_schedule_bits_d_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_schedule_bits_d_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_schedule_bits_d_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [11:0] abc_mshrs_2_io_schedule_bits_d_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [5:0] abc_mshrs_2_io_schedule_bits_d_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [5:0] abc_mshrs_2_io_schedule_bits_d_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [9:0] abc_mshrs_2_io_schedule_bits_d_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_schedule_bits_d_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_d_bits_bad; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_e_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_schedule_bits_e_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_x_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_dir_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [9:0] abc_mshrs_2_io_schedule_bits_dir_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_schedule_bits_dir_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [1:0] abc_mshrs_2_io_schedule_bits_dir_bits_data_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_dir_bits_data_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [11:0] abc_mshrs_2_io_schedule_bits_dir_bits_data_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_schedule_bits_reload; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_sinkc_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_sinkc_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [11:0] abc_mshrs_2_io_sinkc_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_sinkc_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_sinkc_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_sinkc_bits_data; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_sinkd_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_sinkd_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_sinkd_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_sinkd_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [2:0] abc_mshrs_2_io_sinkd_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_sinkd_bits_denied; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_sinke_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [9:0] abc_mshrs_2_io_nestedwb_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire [11:0] abc_mshrs_2_io_nestedwb_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_nestedwb_b_toN; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_nestedwb_b_toB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_nestedwb_b_clr_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_2_io_nestedwb_c_set_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
  wire  abc_mshrs_3_clock; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_reset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_allocate_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_allocate_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_allocate_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_allocate_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_allocate_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_allocate_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_allocate_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_allocate_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_allocate_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [11:0] abc_mshrs_3_io_allocate_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [5:0] abc_mshrs_3_io_allocate_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [5:0] abc_mshrs_3_io_allocate_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [9:0] abc_mshrs_3_io_allocate_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_allocate_bits_repeat; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_directory_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_directory_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [1:0] abc_mshrs_3_io_directory_bits_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_directory_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [11:0] abc_mshrs_3_io_directory_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_directory_bits_hit; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_directory_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_status_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [9:0] abc_mshrs_3_io_status_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [11:0] abc_mshrs_3_io_status_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_status_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_status_bits_blockB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_status_bits_nestB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_status_bits_blockC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_status_bits_nestC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_ready; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_a_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [11:0] abc_mshrs_3_io_schedule_bits_a_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [9:0] abc_mshrs_3_io_schedule_bits_a_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_schedule_bits_a_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_a_bits_block; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_b_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_schedule_bits_b_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [11:0] abc_mshrs_3_io_schedule_bits_b_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [9:0] abc_mshrs_3_io_schedule_bits_b_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_b_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_c_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_schedule_bits_c_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_schedule_bits_c_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [11:0] abc_mshrs_3_io_schedule_bits_c_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [9:0] abc_mshrs_3_io_schedule_bits_c_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_schedule_bits_c_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_c_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_d_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_d_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_d_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_d_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_d_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_schedule_bits_d_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_schedule_bits_d_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_schedule_bits_d_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_schedule_bits_d_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [11:0] abc_mshrs_3_io_schedule_bits_d_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [5:0] abc_mshrs_3_io_schedule_bits_d_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [5:0] abc_mshrs_3_io_schedule_bits_d_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [9:0] abc_mshrs_3_io_schedule_bits_d_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_schedule_bits_d_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_d_bits_bad; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_e_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_schedule_bits_e_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_x_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_dir_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [9:0] abc_mshrs_3_io_schedule_bits_dir_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_schedule_bits_dir_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [1:0] abc_mshrs_3_io_schedule_bits_dir_bits_data_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_dir_bits_data_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [11:0] abc_mshrs_3_io_schedule_bits_dir_bits_data_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_schedule_bits_reload; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_sinkc_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_sinkc_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [11:0] abc_mshrs_3_io_sinkc_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_sinkc_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_sinkc_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_sinkc_bits_data; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_sinkd_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_sinkd_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_sinkd_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_sinkd_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [2:0] abc_mshrs_3_io_sinkd_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_sinkd_bits_denied; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_sinke_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [9:0] abc_mshrs_3_io_nestedwb_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire [11:0] abc_mshrs_3_io_nestedwb_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_nestedwb_b_toN; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_nestedwb_b_toB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_nestedwb_b_clr_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_3_io_nestedwb_c_set_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
  wire  abc_mshrs_4_clock; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_reset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_allocate_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_allocate_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_allocate_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_allocate_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_allocate_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_allocate_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_allocate_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_allocate_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_allocate_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [11:0] abc_mshrs_4_io_allocate_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [5:0] abc_mshrs_4_io_allocate_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [5:0] abc_mshrs_4_io_allocate_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [9:0] abc_mshrs_4_io_allocate_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_allocate_bits_repeat; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_directory_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_directory_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [1:0] abc_mshrs_4_io_directory_bits_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_directory_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [11:0] abc_mshrs_4_io_directory_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_directory_bits_hit; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_directory_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_status_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [9:0] abc_mshrs_4_io_status_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [11:0] abc_mshrs_4_io_status_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_status_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_status_bits_blockB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_status_bits_nestB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_status_bits_blockC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_status_bits_nestC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_ready; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_a_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [11:0] abc_mshrs_4_io_schedule_bits_a_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [9:0] abc_mshrs_4_io_schedule_bits_a_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_schedule_bits_a_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_a_bits_block; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_b_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_schedule_bits_b_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [11:0] abc_mshrs_4_io_schedule_bits_b_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [9:0] abc_mshrs_4_io_schedule_bits_b_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_b_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_c_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_schedule_bits_c_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_schedule_bits_c_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [11:0] abc_mshrs_4_io_schedule_bits_c_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [9:0] abc_mshrs_4_io_schedule_bits_c_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_schedule_bits_c_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_c_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_d_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_d_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_d_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_d_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_d_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_schedule_bits_d_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_schedule_bits_d_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_schedule_bits_d_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_schedule_bits_d_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [11:0] abc_mshrs_4_io_schedule_bits_d_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [5:0] abc_mshrs_4_io_schedule_bits_d_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [5:0] abc_mshrs_4_io_schedule_bits_d_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [9:0] abc_mshrs_4_io_schedule_bits_d_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_schedule_bits_d_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_d_bits_bad; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_e_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_schedule_bits_e_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_x_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_dir_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [9:0] abc_mshrs_4_io_schedule_bits_dir_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_schedule_bits_dir_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [1:0] abc_mshrs_4_io_schedule_bits_dir_bits_data_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_dir_bits_data_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [11:0] abc_mshrs_4_io_schedule_bits_dir_bits_data_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_schedule_bits_reload; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_sinkc_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_sinkc_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [11:0] abc_mshrs_4_io_sinkc_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_sinkc_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_sinkc_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_sinkc_bits_data; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_sinkd_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_sinkd_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_sinkd_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_sinkd_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [2:0] abc_mshrs_4_io_sinkd_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_sinkd_bits_denied; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_sinke_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [9:0] abc_mshrs_4_io_nestedwb_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire [11:0] abc_mshrs_4_io_nestedwb_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_nestedwb_b_toN; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_nestedwb_b_toB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_nestedwb_b_clr_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  abc_mshrs_4_io_nestedwb_c_set_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
  wire  bc_mshr_clock; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_reset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_allocate_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_allocate_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_allocate_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_allocate_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_allocate_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_allocate_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_allocate_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_allocate_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_allocate_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [11:0] bc_mshr_io_allocate_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [5:0] bc_mshr_io_allocate_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [5:0] bc_mshr_io_allocate_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [9:0] bc_mshr_io_allocate_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_allocate_bits_repeat; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_directory_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_directory_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [1:0] bc_mshr_io_directory_bits_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_directory_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [11:0] bc_mshr_io_directory_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_directory_bits_hit; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_directory_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_status_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [9:0] bc_mshr_io_status_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [11:0] bc_mshr_io_status_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_status_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_status_bits_blockB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_status_bits_nestB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_status_bits_blockC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_status_bits_nestC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_ready; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_a_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [11:0] bc_mshr_io_schedule_bits_a_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [9:0] bc_mshr_io_schedule_bits_a_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_schedule_bits_a_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_a_bits_block; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_b_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_schedule_bits_b_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [11:0] bc_mshr_io_schedule_bits_b_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [9:0] bc_mshr_io_schedule_bits_b_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_b_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_c_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_schedule_bits_c_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_schedule_bits_c_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [11:0] bc_mshr_io_schedule_bits_c_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [9:0] bc_mshr_io_schedule_bits_c_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_schedule_bits_c_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_c_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_d_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_d_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_d_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_d_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_d_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_schedule_bits_d_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_schedule_bits_d_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_schedule_bits_d_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_schedule_bits_d_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [11:0] bc_mshr_io_schedule_bits_d_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [5:0] bc_mshr_io_schedule_bits_d_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [5:0] bc_mshr_io_schedule_bits_d_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [9:0] bc_mshr_io_schedule_bits_d_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_schedule_bits_d_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_d_bits_bad; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_e_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_schedule_bits_e_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_x_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_dir_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [9:0] bc_mshr_io_schedule_bits_dir_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_schedule_bits_dir_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [1:0] bc_mshr_io_schedule_bits_dir_bits_data_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_dir_bits_data_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [11:0] bc_mshr_io_schedule_bits_dir_bits_data_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_schedule_bits_reload; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_sinkc_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_sinkc_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [11:0] bc_mshr_io_sinkc_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_sinkc_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_sinkc_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_sinkc_bits_data; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_sinkd_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_sinkd_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_sinkd_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_sinkd_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [2:0] bc_mshr_io_sinkd_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_sinkd_bits_denied; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_sinke_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [9:0] bc_mshr_io_nestedwb_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire [11:0] bc_mshr_io_nestedwb_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_nestedwb_b_toN; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_nestedwb_b_toB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_nestedwb_b_clr_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  bc_mshr_io_nestedwb_c_set_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
  wire  c_mshr_clock; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_reset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_allocate_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_allocate_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_allocate_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_allocate_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_allocate_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_allocate_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_allocate_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_allocate_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_allocate_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [11:0] c_mshr_io_allocate_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [5:0] c_mshr_io_allocate_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [5:0] c_mshr_io_allocate_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [9:0] c_mshr_io_allocate_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_allocate_bits_repeat; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_directory_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_directory_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [1:0] c_mshr_io_directory_bits_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_directory_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [11:0] c_mshr_io_directory_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_directory_bits_hit; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_directory_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_status_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [9:0] c_mshr_io_status_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [11:0] c_mshr_io_status_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_status_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_status_bits_blockB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_status_bits_nestB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_status_bits_blockC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_status_bits_nestC; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_ready; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_a_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [11:0] c_mshr_io_schedule_bits_a_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [9:0] c_mshr_io_schedule_bits_a_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_schedule_bits_a_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_a_bits_block; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_b_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_schedule_bits_b_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [11:0] c_mshr_io_schedule_bits_b_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [9:0] c_mshr_io_schedule_bits_b_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_b_bits_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_c_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_schedule_bits_c_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_schedule_bits_c_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [11:0] c_mshr_io_schedule_bits_c_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [9:0] c_mshr_io_schedule_bits_c_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_schedule_bits_c_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_c_bits_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_d_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_d_bits_prio_0; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_d_bits_prio_1; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_d_bits_prio_2; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_d_bits_control; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_schedule_bits_d_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_schedule_bits_d_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_schedule_bits_d_bits_size; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_schedule_bits_d_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [11:0] c_mshr_io_schedule_bits_d_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [5:0] c_mshr_io_schedule_bits_d_bits_offset; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [5:0] c_mshr_io_schedule_bits_d_bits_put; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [9:0] c_mshr_io_schedule_bits_d_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_schedule_bits_d_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_d_bits_bad; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_e_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_schedule_bits_e_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_x_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_dir_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [9:0] c_mshr_io_schedule_bits_dir_bits_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_schedule_bits_dir_bits_way; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [1:0] c_mshr_io_schedule_bits_dir_bits_data_state; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_dir_bits_data_clients; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [11:0] c_mshr_io_schedule_bits_dir_bits_data_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_schedule_bits_reload; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_sinkc_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_sinkc_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [11:0] c_mshr_io_sinkc_bits_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_sinkc_bits_source; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_sinkc_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_sinkc_bits_data; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_sinkd_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_sinkd_bits_last; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_sinkd_bits_opcode; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_sinkd_bits_param; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [2:0] c_mshr_io_sinkd_bits_sink; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_sinkd_bits_denied; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_sinke_valid; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [9:0] c_mshr_io_nestedwb_set; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire [11:0] c_mshr_io_nestedwb_tag; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_nestedwb_b_toN; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_nestedwb_b_toB; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_nestedwb_b_clr_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  c_mshr_io_nestedwb_c_set_dirty; // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
  wire  _T; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100127.4]
  wire  _T_2; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100130.4]
  wire  _T_4; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100133.4]
  wire  _T_6; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100140.4]
  wire  _T_8; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100143.4]
  wire  _T_10; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100146.4]
  wire  _T_12; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100153.4]
  wire  _T_14; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100156.4]
  wire  _T_16; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100159.4]
  wire  _T_18; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100166.4]
  wire  _T_20; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100169.4]
  wire  _T_22; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100172.4]
  wire  _T_24; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100179.4]
  wire  _T_26; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100182.4]
  wire  _T_28; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100185.4]
  wire  _T_30; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100192.4]
  wire  _T_32; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100195.4]
  wire  _T_34; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100198.4]
  wire  _T_36; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100205.4]
  wire  _T_38; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100208.4]
  wire  _T_40; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100211.4]
  wire  _T_42; // @[Scheduler.scala 88:54:chipyard.TestHarness.RocketConfig.fir@100218.4]
  wire  _T_43; // @[Scheduler.scala 88:30:chipyard.TestHarness.RocketConfig.fir@100219.4]
  wire  _T_44; // @[Scheduler.scala 89:54:chipyard.TestHarness.RocketConfig.fir@100220.4]
  wire  _T_45; // @[Scheduler.scala 89:30:chipyard.TestHarness.RocketConfig.fir@100221.4]
  wire  mshr_stall_0; // @[Scheduler.scala 88:86:chipyard.TestHarness.RocketConfig.fir@100222.4]
  wire  _T_46; // @[Scheduler.scala 88:54:chipyard.TestHarness.RocketConfig.fir@100223.4]
  wire  _T_47; // @[Scheduler.scala 88:30:chipyard.TestHarness.RocketConfig.fir@100224.4]
  wire  _T_48; // @[Scheduler.scala 89:54:chipyard.TestHarness.RocketConfig.fir@100225.4]
  wire  _T_49; // @[Scheduler.scala 89:30:chipyard.TestHarness.RocketConfig.fir@100226.4]
  wire  mshr_stall_1; // @[Scheduler.scala 88:86:chipyard.TestHarness.RocketConfig.fir@100227.4]
  wire  _T_50; // @[Scheduler.scala 88:54:chipyard.TestHarness.RocketConfig.fir@100228.4]
  wire  _T_51; // @[Scheduler.scala 88:30:chipyard.TestHarness.RocketConfig.fir@100229.4]
  wire  _T_52; // @[Scheduler.scala 89:54:chipyard.TestHarness.RocketConfig.fir@100230.4]
  wire  _T_53; // @[Scheduler.scala 89:30:chipyard.TestHarness.RocketConfig.fir@100231.4]
  wire  mshr_stall_2; // @[Scheduler.scala 88:86:chipyard.TestHarness.RocketConfig.fir@100232.4]
  wire  _T_54; // @[Scheduler.scala 88:54:chipyard.TestHarness.RocketConfig.fir@100233.4]
  wire  _T_55; // @[Scheduler.scala 88:30:chipyard.TestHarness.RocketConfig.fir@100234.4]
  wire  _T_56; // @[Scheduler.scala 89:54:chipyard.TestHarness.RocketConfig.fir@100235.4]
  wire  _T_57; // @[Scheduler.scala 89:30:chipyard.TestHarness.RocketConfig.fir@100236.4]
  wire  mshr_stall_3; // @[Scheduler.scala 88:86:chipyard.TestHarness.RocketConfig.fir@100237.4]
  wire  _T_58; // @[Scheduler.scala 88:54:chipyard.TestHarness.RocketConfig.fir@100238.4]
  wire  _T_59; // @[Scheduler.scala 88:30:chipyard.TestHarness.RocketConfig.fir@100239.4]
  wire  _T_60; // @[Scheduler.scala 89:54:chipyard.TestHarness.RocketConfig.fir@100240.4]
  wire  _T_61; // @[Scheduler.scala 89:30:chipyard.TestHarness.RocketConfig.fir@100241.4]
  wire  mshr_stall_4; // @[Scheduler.scala 88:86:chipyard.TestHarness.RocketConfig.fir@100242.4]
  wire  _T_62; // @[Scheduler.scala 92:58:chipyard.TestHarness.RocketConfig.fir@100243.4]
  wire  mshr_stall_5; // @[Scheduler.scala 92:28:chipyard.TestHarness.RocketConfig.fir@100244.4]
  wire  _T_67; // @[Scheduler.scala 105:28:chipyard.TestHarness.RocketConfig.fir@100254.4]
  wire  _T_68; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100255.4]
  wire  _T_69; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100256.4]
  wire  _T_70; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100257.4]
  wire  _T_71; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100258.4]
  wire  _T_72; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100259.4]
  wire  _T_73; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100260.4]
  wire  _T_74; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100261.4]
  wire  _T_75; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100262.4]
  wire  _T_76; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100263.4]
  wire  _T_77; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100264.4]
  wire  _T_78; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100265.4]
  wire  _T_79; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100266.4]
  wire  _T_80; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100267.4]
  wire  _T_81; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100268.4]
  wire  _T_82; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100269.4]
  wire  _T_83; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100270.4]
  wire  _T_84; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100271.4]
  wire  _T_85; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100272.4]
  wire  _T_86; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100273.4]
  wire  _T_87; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100274.4]
  wire  _T_88; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100275.4]
  wire  _T_89; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100276.4]
  wire  _T_90; // @[Scheduler.scala 105:28:chipyard.TestHarness.RocketConfig.fir@100277.4]
  wire  _T_91; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100278.4]
  wire  _T_92; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100279.4]
  wire  _T_93; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100280.4]
  wire  _T_94; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100281.4]
  wire  _T_95; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100282.4]
  wire  _T_96; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100283.4]
  wire  _T_97; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100284.4]
  wire  _T_98; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100285.4]
  wire  _T_99; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100286.4]
  wire  _T_100; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100287.4]
  wire  _T_101; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100288.4]
  wire  _T_102; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100289.4]
  wire  _T_103; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100290.4]
  wire  _T_104; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100291.4]
  wire  _T_105; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100292.4]
  wire  _T_106; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100293.4]
  wire  _T_107; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100294.4]
  wire  _T_108; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100295.4]
  wire  _T_109; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100296.4]
  wire  _T_110; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100297.4]
  wire  _T_111; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100298.4]
  wire  _T_112; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100299.4]
  wire  _T_113; // @[Scheduler.scala 105:28:chipyard.TestHarness.RocketConfig.fir@100300.4]
  wire  _T_114; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100301.4]
  wire  _T_115; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100302.4]
  wire  _T_116; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100303.4]
  wire  _T_117; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100304.4]
  wire  _T_118; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100305.4]
  wire  _T_119; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100306.4]
  wire  _T_120; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100307.4]
  wire  _T_121; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100308.4]
  wire  _T_122; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100309.4]
  wire  _T_123; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100310.4]
  wire  _T_124; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100311.4]
  wire  _T_125; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100312.4]
  wire  _T_126; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100313.4]
  wire  _T_127; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100314.4]
  wire  _T_128; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100315.4]
  wire  _T_129; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100316.4]
  wire  _T_130; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100317.4]
  wire  _T_131; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100318.4]
  wire  _T_132; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100319.4]
  wire  _T_133; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100320.4]
  wire  _T_134; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100321.4]
  wire  _T_135; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100322.4]
  wire  _T_136; // @[Scheduler.scala 105:28:chipyard.TestHarness.RocketConfig.fir@100323.4]
  wire  _T_137; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100324.4]
  wire  _T_138; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100325.4]
  wire  _T_139; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100326.4]
  wire  _T_140; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100327.4]
  wire  _T_141; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100328.4]
  wire  _T_142; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100329.4]
  wire  _T_143; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100330.4]
  wire  _T_144; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100331.4]
  wire  _T_145; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100332.4]
  wire  _T_146; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100333.4]
  wire  _T_147; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100334.4]
  wire  _T_148; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100335.4]
  wire  _T_149; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100336.4]
  wire  _T_150; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100337.4]
  wire  _T_151; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100338.4]
  wire  _T_152; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100339.4]
  wire  _T_153; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100340.4]
  wire  _T_154; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100341.4]
  wire  _T_155; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100342.4]
  wire  _T_156; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100343.4]
  wire  _T_157; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100344.4]
  wire  _T_158; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100345.4]
  wire  _T_159; // @[Scheduler.scala 105:28:chipyard.TestHarness.RocketConfig.fir@100346.4]
  wire  _T_160; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100347.4]
  wire  _T_161; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100348.4]
  wire  _T_162; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100349.4]
  wire  _T_163; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100350.4]
  wire  _T_164; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100351.4]
  wire  _T_165; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100352.4]
  wire  _T_166; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100353.4]
  wire  _T_167; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100354.4]
  wire  _T_168; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100355.4]
  wire  _T_169; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100356.4]
  wire  _T_170; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100357.4]
  wire  _T_171; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100358.4]
  wire  _T_172; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100359.4]
  wire  _T_173; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100360.4]
  wire  _T_174; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100361.4]
  wire  _T_175; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100362.4]
  wire  _T_176; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100363.4]
  wire  _T_177; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100364.4]
  wire  _T_178; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100365.4]
  wire  _T_179; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100366.4]
  wire  _T_180; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100367.4]
  wire  _T_181; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100368.4]
  wire  _T_182; // @[Scheduler.scala 105:28:chipyard.TestHarness.RocketConfig.fir@100369.4]
  wire  _T_183; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100370.4]
  wire  _T_184; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100371.4]
  wire  _T_185; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100372.4]
  wire  _T_186; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100373.4]
  wire  _T_187; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100374.4]
  wire  _T_188; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100375.4]
  wire  _T_189; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100376.4]
  wire  _T_190; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100377.4]
  wire  _T_191; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100378.4]
  wire  _T_192; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100379.4]
  wire  _T_193; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100380.4]
  wire  _T_194; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100381.4]
  wire  _T_195; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100382.4]
  wire  _T_196; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100383.4]
  wire  _T_197; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100384.4]
  wire  _T_198; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100385.4]
  wire  _T_199; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100386.4]
  wire  _T_200; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100387.4]
  wire  _T_201; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100388.4]
  wire  _T_202; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100389.4]
  wire  _T_203; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100390.4]
  wire  _T_204; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100391.4]
  wire  _T_206; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100393.4]
  wire  _T_207; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100394.4]
  wire  _T_208; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100395.4]
  wire  _T_209; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100396.4]
  wire  _T_210; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100397.4]
  wire  _T_211; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100398.4]
  wire  _T_212; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100399.4]
  wire  _T_213; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100400.4]
  wire  _T_214; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100401.4]
  wire  _T_215; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100402.4]
  wire  _T_216; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100403.4]
  wire  _T_217; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100404.4]
  wire  _T_218; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100405.4]
  wire  _T_219; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100406.4]
  wire  _T_220; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100407.4]
  wire  _T_221; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100408.4]
  wire  _T_222; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100409.4]
  wire  _T_223; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100410.4]
  wire  _T_224; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100411.4]
  wire  _T_225; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100412.4]
  wire  _T_226; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100413.4]
  wire  _T_227; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100414.4]
  wire [6:0] mshr_request; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@100420.4]
  reg [6:0] robin_filter; // @[Scheduler.scala 116:29:chipyard.TestHarness.RocketConfig.fir@100421.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_233; // @[Scheduler.scala 117:54:chipyard.TestHarness.RocketConfig.fir@100422.4]
  wire [13:0] robin_request; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@100423.4]
  wire [14:0] _T_234; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@100424.4]
  wire [13:0] _T_236; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@100426.4]
  wire [15:0] _T_237; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@100427.4]
  wire [13:0] _T_239; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@100429.4]
  wire [17:0] _T_240; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@100430.4]
  wire [13:0] _T_242; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@100432.4]
  wire [21:0] _T_243; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@100433.4]
  wire [13:0] _T_245; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@100435.4]
  wire [14:0] _T_247; // @[Scheduler.scala 118:48:chipyard.TestHarness.RocketConfig.fir@100437.4]
  wire [14:0] _T_248; // @[Scheduler.scala 118:24:chipyard.TestHarness.RocketConfig.fir@100438.4]
  wire [14:0] _GEN_141; // @[Scheduler.scala 118:54:chipyard.TestHarness.RocketConfig.fir@100439.4]
  wire [14:0] mshr_selectOH2; // @[Scheduler.scala 118:54:chipyard.TestHarness.RocketConfig.fir@100439.4]
  wire [6:0] mshr_selectOH; // @[Scheduler.scala 119:70:chipyard.TestHarness.RocketConfig.fir@100442.4]
  wire  _T_253; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@100445.4]
  wire [3:0] _GEN_142; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@100446.4]
  wire [3:0] _T_254; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@100446.4]
  wire  _T_257; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@100449.4]
  wire [1:0] _T_258; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@100450.4]
  wire [1:0] _T_260; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@100452.4]
  wire [2:0] mshr_select; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@100453.4]
  wire [16:0] _T_271; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100464.4]
  wire [35:0] _T_277; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100470.4]
  wire [23:0] _T_282; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100475.4]
  wire [89:0] _T_289; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100482.4]
  wire [5:0] _T_294; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100487.4]
  wire [39:0] _T_300; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100493.4]
  wire [27:0] _T_305; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100498.4]
  wire [187:0] _T_313; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100506.4]
  wire [187:0] _T_314; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100507.4]
  wire [16:0] _T_318; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100511.4]
  wire [35:0] _T_324; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100517.4]
  wire [23:0] _T_329; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100522.4]
  wire [89:0] _T_336; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100529.4]
  wire [5:0] _T_341; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100534.4]
  wire [39:0] _T_347; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100540.4]
  wire [27:0] _T_352; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100545.4]
  wire [187:0] _T_360; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100553.4]
  wire [187:0] _T_361; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100554.4]
  wire [16:0] _T_365; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100558.4]
  wire [35:0] _T_371; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100564.4]
  wire [23:0] _T_376; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100569.4]
  wire [89:0] _T_383; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100576.4]
  wire [5:0] _T_388; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100581.4]
  wire [39:0] _T_394; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100587.4]
  wire [27:0] _T_399; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100592.4]
  wire [187:0] _T_407; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100600.4]
  wire [187:0] _T_408; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100601.4]
  wire [16:0] _T_412; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100605.4]
  wire [35:0] _T_418; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100611.4]
  wire [23:0] _T_423; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100616.4]
  wire [89:0] _T_430; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100623.4]
  wire [5:0] _T_435; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100628.4]
  wire [39:0] _T_441; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100634.4]
  wire [27:0] _T_446; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100639.4]
  wire [187:0] _T_454; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100647.4]
  wire [187:0] _T_455; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100648.4]
  wire [16:0] _T_459; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100652.4]
  wire [35:0] _T_465; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100658.4]
  wire [23:0] _T_470; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100663.4]
  wire [89:0] _T_477; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100670.4]
  wire [5:0] _T_482; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100675.4]
  wire [39:0] _T_488; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100681.4]
  wire [27:0] _T_493; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100686.4]
  wire [187:0] _T_501; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100694.4]
  wire [187:0] _T_502; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100695.4]
  wire [16:0] _T_506; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100699.4]
  wire [35:0] _T_512; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100705.4]
  wire [23:0] _T_517; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100710.4]
  wire [89:0] _T_524; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100717.4]
  wire [5:0] _T_529; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100722.4]
  wire [39:0] _T_535; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100728.4]
  wire [27:0] _T_540; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100733.4]
  wire [187:0] _T_548; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100741.4]
  wire [187:0] _T_549; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100742.4]
  wire [16:0] _T_553; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100746.4]
  wire [35:0] _T_559; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100752.4]
  wire [23:0] _T_564; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100757.4]
  wire [89:0] _T_571; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100764.4]
  wire [5:0] _T_576; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100769.4]
  wire [39:0] _T_582; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100775.4]
  wire [27:0] _T_587; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100780.4]
  wire [187:0] _T_595; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100788.4]
  wire [187:0] _T_596; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100789.4]
  wire [187:0] _T_597; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100790.4]
  wire [187:0] _T_598; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100791.4]
  wire [187:0] _T_599; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100792.4]
  wire [187:0] _T_600; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100793.4]
  wire [187:0] _T_601; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100794.4]
  wire [187:0] _T_602; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100795.4]
  wire  schedule_reload; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100799.4]
  wire [2:0] schedule_c_bits_opcode; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100867.4]
  wire [11:0] _T_658; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100900.4]
  wire [11:0] _T_659; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100901.4]
  wire [11:0] _T_660; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100902.4]
  wire [11:0] _T_661; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100903.4]
  wire [11:0] _T_662; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100904.4]
  wire [11:0] _T_663; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100905.4]
  wire [11:0] _T_664; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100906.4]
  wire [11:0] _T_665; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100907.4]
  wire [11:0] _T_666; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100908.4]
  wire [11:0] _T_667; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100909.4]
  wire [11:0] _T_668; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100910.4]
  wire [11:0] _T_669; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100911.4]
  wire [11:0] scheduleTag; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100912.4]
  wire [9:0] _T_678; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100922.4]
  wire [9:0] _T_679; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100923.4]
  wire [9:0] _T_680; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100924.4]
  wire [9:0] _T_681; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100925.4]
  wire [9:0] _T_682; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100926.4]
  wire [9:0] _T_683; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100927.4]
  wire [9:0] _T_684; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100928.4]
  wire [9:0] _T_685; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100929.4]
  wire [9:0] _T_686; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100930.4]
  wire [9:0] _T_687; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100931.4]
  wire [9:0] _T_688; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100932.4]
  wire [9:0] _T_689; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100933.4]
  wire [9:0] scheduleSet; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100934.4]
  wire  _T_691; // @[Scheduler.scala 126:25:chipyard.TestHarness.RocketConfig.fir@100937.4]
  wire [6:0] _GEN_143; // @[package.scala 208:43:chipyard.TestHarness.RocketConfig.fir@100940.6]
  wire [6:0] _T_693; // @[package.scala 208:43:chipyard.TestHarness.RocketConfig.fir@100940.6]
  wire [6:0] _GEN_144; // @[package.scala 208:43:chipyard.TestHarness.RocketConfig.fir@100942.6]
  wire [6:0] _T_695; // @[package.scala 208:43:chipyard.TestHarness.RocketConfig.fir@100942.6]
  wire [6:0] _GEN_145; // @[package.scala 208:43:chipyard.TestHarness.RocketConfig.fir@100944.6]
  wire [6:0] _T_697; // @[package.scala 208:43:chipyard.TestHarness.RocketConfig.fir@100944.6]
  wire [6:0] _T_699; // @[Scheduler.scala 126:47:chipyard.TestHarness.RocketConfig.fir@100946.6]
  wire  _T_704; // @[Scheduler.scala 146:37:chipyard.TestHarness.RocketConfig.fir@100967.4]
  wire  _T_705; // @[Scheduler.scala 146:123:chipyard.TestHarness.RocketConfig.fir@100968.4]
  wire  _T_708; // @[Scheduler.scala 147:123:chipyard.TestHarness.RocketConfig.fir@100972.4]
  wire  _T_711; // @[Scheduler.scala 149:37:chipyard.TestHarness.RocketConfig.fir@100977.4]
  wire  _T_713; // @[Scheduler.scala 153:62:chipyard.TestHarness.RocketConfig.fir@100982.4]
  wire  _T_714; // @[Scheduler.scala 153:84:chipyard.TestHarness.RocketConfig.fir@100983.4]
  wire  request_valid; // @[Scheduler.scala 153:39:chipyard.TestHarness.RocketConfig.fir@100984.4]
  wire  _T_716_control; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  wire [2:0] _T_716_opcode; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  wire [2:0] _T_716_param; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  wire [2:0] _T_716_size; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  wire [2:0] _T_716_source; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  wire [11:0] _T_716_tag; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  wire [5:0] _T_716_offset; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  wire [5:0] _T_716_put; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  wire [9:0] _T_716_set; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  wire  request_bits_prio_0; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  wire  request_bits_prio_2; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  wire  request_bits_control; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  wire [2:0] request_bits_opcode; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  wire [2:0] request_bits_param; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  wire [2:0] request_bits_size; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  wire [2:0] request_bits_source; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  wire [11:0] request_bits_tag; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  wire [5:0] request_bits_offset; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  wire [5:0] request_bits_put; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  wire [9:0] request_bits_set; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  wire  _T_739; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101013.4]
  wire  _T_740; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101014.4]
  wire  _T_737; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101011.4]
  wire  _T_738; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101012.4]
  wire  _T_735; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101009.4]
  wire  _T_736; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101010.4]
  wire  _T_733; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101007.4]
  wire  _T_734; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101008.4]
  wire  _T_731; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101005.4]
  wire  _T_732; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101006.4]
  wire  _T_729; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101003.4]
  wire  _T_730; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101004.4]
  wire  _T_727; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101001.4]
  wire  _T_728; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101002.4]
  wire [6:0] setMatches; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101020.4]
  wire  _T_746; // @[Scheduler.scala 162:30:chipyard.TestHarness.RocketConfig.fir@101021.4]
  wire  alloc; // @[Scheduler.scala 162:15:chipyard.TestHarness.RocketConfig.fir@101022.4]
  wire [20:0] _T_849; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101137.4]
  wire [20:0] selected_requests; // @[Scheduler.scala 195:76:chipyard.TestHarness.RocketConfig.fir@101138.4]
  wire  a_pop; // @[Scheduler.scala 196:82:chipyard.TestHarness.RocketConfig.fir@101140.4]
  wire  b_pop; // @[Scheduler.scala 197:82:chipyard.TestHarness.RocketConfig.fir@101142.4]
  wire  _T_862; // @[Scheduler.scala 201:23:chipyard.TestHarness.RocketConfig.fir@101155.4]
  wire  c_pop; // @[Scheduler.scala 198:82:chipyard.TestHarness.RocketConfig.fir@101144.4]
  wire  may_pop; // @[Scheduler.scala 201:32:chipyard.TestHarness.RocketConfig.fir@101156.4]
  wire  _T_1062; // @[Scheduler.scala 236:64:chipyard.TestHarness.RocketConfig.fir@101413.4]
  wire  lb_tag_mismatch; // @[Scheduler.scala 235:37:chipyard.TestHarness.RocketConfig.fir@101412.4]
  wire  mshr_uses_directory_assuming_no_bypass; // @[Scheduler.scala 236:75:chipyard.TestHarness.RocketConfig.fir@101414.4]
  wire  _T_1072; // @[Scheduler.scala 247:16:chipyard.TestHarness.RocketConfig.fir@101429.4]
  wire  _T_1073; // @[Scheduler.scala 247:13:chipyard.TestHarness.RocketConfig.fir@101430.4]
  wire [6:0] mshr_validOH; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101424.4]
  wire [6:0] _T_1070; // @[Scheduler.scala 242:20:chipyard.TestHarness.RocketConfig.fir@101425.4]
  wire  _T_831; // @[Scheduler.scala 171:46:chipyard.TestHarness.RocketConfig.fir@101115.4]
  wire [6:0] prioFilter; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101118.4]
  wire [6:0] _T_1071; // @[Scheduler.scala 242:34:chipyard.TestHarness.RocketConfig.fir@101426.4]
  wire  mshr_free; // @[Scheduler.scala 242:51:chipyard.TestHarness.RocketConfig.fir@101427.4]
  wire  _T_1074; // @[Scheduler.scala 247:56:chipyard.TestHarness.RocketConfig.fir@101431.4]
  wire  _T_1079; // @[Scheduler.scala 248:87:chipyard.TestHarness.RocketConfig.fir@101436.4]
  wire  _T_817; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101099.4]
  wire  _T_818; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101100.4]
  wire  _T_824; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101106.4]
  wire  _T_819; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101101.4]
  wire  _T_825; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101107.4]
  wire  _T_820; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101102.4]
  wire  _T_826; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101108.4]
  wire  _T_821; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101103.4]
  wire  _T_827; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101109.4]
  wire  _T_822; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101104.4]
  wire  _T_828; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101110.4]
  wire  _T_823; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101105.4]
  wire  _T_829; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101111.4]
  wire  nestC; // @[Scheduler.scala 169:70:chipyard.TestHarness.RocketConfig.fir@101114.4]
  wire  _T_1083; // @[Scheduler.scala 249:13:chipyard.TestHarness.RocketConfig.fir@101440.4]
  wire  _T_1085; // @[Scheduler.scala 249:56:chipyard.TestHarness.RocketConfig.fir@101442.4]
  wire  request_alloc_cases; // @[Scheduler.scala 248:112:chipyard.TestHarness.RocketConfig.fir@101443.4]
  wire [6:0] lowerMatches; // @[Scheduler.scala 172:33:chipyard.TestHarness.RocketConfig.fir@101119.4]
  wire  _T_834; // @[Scheduler.scala 174:31:chipyard.TestHarness.RocketConfig.fir@101120.4]
  wire  _T_837; // @[Scheduler.scala 174:47:chipyard.TestHarness.RocketConfig.fir@101123.4]
  wire  _T_838; // @[Scheduler.scala 174:44:chipyard.TestHarness.RocketConfig.fir@101124.4]
  wire  _T_775; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101053.4]
  wire  _T_776; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101054.4]
  wire  _T_782; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101060.4]
  wire  _T_777; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101055.4]
  wire  _T_783; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101061.4]
  wire  _T_778; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101056.4]
  wire  _T_784; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101062.4]
  wire  _T_779; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101057.4]
  wire  _T_785; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101063.4]
  wire  _T_780; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101058.4]
  wire  _T_786; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101064.4]
  wire  _T_781; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101059.4]
  wire  _T_787; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101065.4]
  wire  blockC; // @[Scheduler.scala 165:70:chipyard.TestHarness.RocketConfig.fir@101068.4]
  wire  _T_841; // @[Scheduler.scala 174:68:chipyard.TestHarness.RocketConfig.fir@101127.4]
  wire  queue; // @[Scheduler.scala 174:65:chipyard.TestHarness.RocketConfig.fir@101128.4]
  wire [6:0] _T_847; // @[Scheduler.scala 190:8:chipyard.TestHarness.RocketConfig.fir@101134.4]
  wire [6:0] lowerMatches1; // @[Scheduler.scala 189:8:chipyard.TestHarness.RocketConfig.fir@101135.4]
  wire [6:0] _T_853; // @[Scheduler.scala 199:38:chipyard.TestHarness.RocketConfig.fir@101145.4]
  wire  _T_854; // @[Scheduler.scala 199:58:chipyard.TestHarness.RocketConfig.fir@101146.4]
  wire  _T_855; // @[Scheduler.scala 200:33:chipyard.TestHarness.RocketConfig.fir@101147.4]
  wire  _T_856; // @[Scheduler.scala 200:58:chipyard.TestHarness.RocketConfig.fir@101148.4]
  wire  _T_858; // @[Scheduler.scala 200:101:chipyard.TestHarness.RocketConfig.fir@101150.4]
  wire  _T_859; // @[Scheduler.scala 200:109:chipyard.TestHarness.RocketConfig.fir@101151.4]
  wire  _T_860; // @[Scheduler.scala 200:69:chipyard.TestHarness.RocketConfig.fir@101152.4]
  wire  _T_861; // @[Scheduler.scala 200:26:chipyard.TestHarness.RocketConfig.fir@101153.4]
  wire  bypassMatches; // @[Scheduler.scala 199:61:chipyard.TestHarness.RocketConfig.fir@101154.4]
  wire  bypassQueue; // @[Scheduler.scala 245:37:chipyard.TestHarness.RocketConfig.fir@101428.4]
  wire  _T_1086; // @[Scheduler.scala 250:66:chipyard.TestHarness.RocketConfig.fir@101444.4]
  wire  _T_1087; // @[Scheduler.scala 250:50:chipyard.TestHarness.RocketConfig.fir@101445.4]
  wire  request_ready; // @[Scheduler.scala 250:40:chipyard.TestHarness.RocketConfig.fir@101446.4]
  wire  _T_718; // @[Scheduler.scala 156:44:chipyard.TestHarness.RocketConfig.fir@100989.4]
  wire  _T_720; // @[Scheduler.scala 157:64:chipyard.TestHarness.RocketConfig.fir@100992.4]
  wire  _T_721; // @[Scheduler.scala 157:61:chipyard.TestHarness.RocketConfig.fir@100993.4]
  wire  _T_725; // @[Scheduler.scala 158:87:chipyard.TestHarness.RocketConfig.fir@100998.4]
  wire  _T_843; // @[Scheduler.scala 182:33:chipyard.TestHarness.RocketConfig.fir@101130.4]
  wire  _T_844; // @[Scheduler.scala 184:31:chipyard.TestHarness.RocketConfig.fir@101131.4]
  wire  bypass; // @[Scheduler.scala 202:39:chipyard.TestHarness.RocketConfig.fir@101158.4]
  wire  _T_864; // @[Scheduler.scala 203:49:chipyard.TestHarness.RocketConfig.fir@101159.4]
  wire  will_reload; // @[Scheduler.scala 203:37:chipyard.TestHarness.RocketConfig.fir@101160.4]
  wire  _T_866; // @[Scheduler.scala 204:48:chipyard.TestHarness.RocketConfig.fir@101162.4]
  wire  will_pop; // @[Scheduler.scala 204:45:chipyard.TestHarness.RocketConfig.fir@101163.4]
  wire  _T_878; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101176.4]
  wire  _T_879; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101177.4]
  wire  _T_881; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101179.4]
  wire  _T_882; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101180.4]
  wire  _T_883; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101181.4]
  wire  _T_884; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101182.4]
  wire  _T_885; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101183.4]
  wire  _T_886; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101184.4]
  wire  _T_887; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101185.4]
  wire  _T_889; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101187.4]
  wire  _T_890; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101188.4]
  wire  _T_891; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101189.4]
  wire  _T_893_prio_0; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  wire  _T_893_prio_1; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  wire  _T_893_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  wire  _T_893_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  wire [2:0] _T_893_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  wire [2:0] _T_893_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  wire [2:0] _T_893_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  wire [2:0] _T_893_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  wire [11:0] _T_893_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  wire [5:0] _T_893_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  wire [5:0] _T_893_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  wire  _T_894; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101196.4]
  wire  _T_895; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101198.4]
  wire  _T_901; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101206.4]
  wire  _T_902; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101207.4]
  wire  _T_904; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101209.4]
  wire  _T_905; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101210.4]
  wire  _T_906; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101211.4]
  wire  _T_907; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101212.4]
  wire  _T_908; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101213.4]
  wire  _T_909; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101214.4]
  wire  _T_910; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101215.4]
  wire  _T_912; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101217.4]
  wire  _T_913; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101218.4]
  wire  _T_914; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101219.4]
  wire  _T_916_prio_0; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  wire  _T_916_prio_1; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  wire  _T_916_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  wire  _T_916_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  wire [2:0] _T_916_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  wire [2:0] _T_916_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  wire [2:0] _T_916_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  wire [2:0] _T_916_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  wire [11:0] _T_916_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  wire [5:0] _T_916_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  wire [5:0] _T_916_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  wire  _T_917; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101226.4]
  wire  _T_918; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101228.4]
  wire  _T_924; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101236.4]
  wire  _T_925; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101237.4]
  wire  _T_927; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101239.4]
  wire  _T_928; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101240.4]
  wire  _T_929; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101241.4]
  wire  _T_930; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101242.4]
  wire  _T_931; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101243.4]
  wire  _T_932; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101244.4]
  wire  _T_933; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101245.4]
  wire  _T_935; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101247.4]
  wire  _T_936; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101248.4]
  wire  _T_937; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101249.4]
  wire  _T_939_prio_0; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  wire  _T_939_prio_1; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  wire  _T_939_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  wire  _T_939_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  wire [2:0] _T_939_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  wire [2:0] _T_939_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  wire [2:0] _T_939_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  wire [2:0] _T_939_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  wire [11:0] _T_939_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  wire [5:0] _T_939_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  wire [5:0] _T_939_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  wire  _T_940; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101256.4]
  wire  _T_941; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101258.4]
  wire  _T_947; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101266.4]
  wire  _T_948; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101267.4]
  wire  _T_950; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101269.4]
  wire  _T_951; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101270.4]
  wire  _T_952; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101271.4]
  wire  _T_953; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101272.4]
  wire  _T_954; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101273.4]
  wire  _T_955; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101274.4]
  wire  _T_956; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101275.4]
  wire  _T_958; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101277.4]
  wire  _T_959; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101278.4]
  wire  _T_960; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101279.4]
  wire  _T_962_prio_0; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  wire  _T_962_prio_1; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  wire  _T_962_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  wire  _T_962_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  wire [2:0] _T_962_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  wire [2:0] _T_962_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  wire [2:0] _T_962_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  wire [2:0] _T_962_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  wire [11:0] _T_962_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  wire [5:0] _T_962_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  wire [5:0] _T_962_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  wire  _T_963; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101286.4]
  wire  _T_964; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101288.4]
  wire  _T_970; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101296.4]
  wire  _T_971; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101297.4]
  wire  _T_973; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101299.4]
  wire  _T_974; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101300.4]
  wire  _T_975; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101301.4]
  wire  _T_976; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101302.4]
  wire  _T_977; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101303.4]
  wire  _T_978; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101304.4]
  wire  _T_979; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101305.4]
  wire  _T_981; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101307.4]
  wire  _T_982; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101308.4]
  wire  _T_983; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101309.4]
  wire  _T_985_prio_0; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  wire  _T_985_prio_1; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  wire  _T_985_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  wire  _T_985_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  wire [2:0] _T_985_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  wire [2:0] _T_985_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  wire [2:0] _T_985_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  wire [2:0] _T_985_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  wire [11:0] _T_985_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  wire [5:0] _T_985_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  wire [5:0] _T_985_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  wire  _T_986; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101316.4]
  wire  _T_987; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101318.4]
  wire  _T_993; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101326.4]
  wire  _T_994; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101327.4]
  wire  _T_996; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101329.4]
  wire  _T_997; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101330.4]
  wire  _T_998; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101331.4]
  wire  _T_999; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101332.4]
  wire  _T_1000; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101333.4]
  wire  _T_1001; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101334.4]
  wire  _T_1002; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101335.4]
  wire  _T_1004; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101337.4]
  wire  _T_1005; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101338.4]
  wire  _T_1006; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101339.4]
  wire  _T_1008_prio_1; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  wire  _T_1008_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  wire  _T_1008_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  wire [2:0] _T_1008_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  wire [2:0] _T_1008_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  wire [2:0] _T_1008_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  wire [2:0] _T_1008_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  wire [11:0] _T_1008_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  wire [5:0] _T_1008_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  wire [5:0] _T_1008_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  wire  _T_1009; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101346.4]
  wire  _T_1010; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101348.4]
  wire  _T_1016; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101356.4]
  wire  _T_1017; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101357.4]
  wire  _T_1019; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101359.4]
  wire  _T_1020; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101360.4]
  wire  _T_1021; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101361.4]
  wire  _T_1022; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101362.4]
  wire  _T_1023; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101363.4]
  wire  _T_1024; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101364.4]
  wire  _T_1025; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101365.4]
  wire  _T_1027; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101367.4]
  wire  _T_1028; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101368.4]
  wire  _T_1029; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101369.4]
  wire  _T_1031_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  wire  _T_1031_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  wire [2:0] _T_1031_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  wire [2:0] _T_1031_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  wire [2:0] _T_1031_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  wire [2:0] _T_1031_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  wire [11:0] _T_1031_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  wire [5:0] _T_1031_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  wire [5:0] _T_1031_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  wire  _T_1032; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101376.4]
  wire  _T_1033; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101378.4]
  wire [20:0] _T_1034; // @[Scheduler.scala 229:25:chipyard.TestHarness.RocketConfig.fir@101380.4]
  wire [20:0] _GEN_146; // @[Scheduler.scala 229:44:chipyard.TestHarness.RocketConfig.fir@101382.4]
  wire [20:0] _T_1036; // @[Scheduler.scala 229:44:chipyard.TestHarness.RocketConfig.fir@101382.4]
  wire [20:0] _GEN_147; // @[Scheduler.scala 229:82:chipyard.TestHarness.RocketConfig.fir@101384.4]
  wire [20:0] _T_1038; // @[Scheduler.scala 229:82:chipyard.TestHarness.RocketConfig.fir@101384.4]
  wire [20:0] prio_requests; // @[Scheduler.scala 229:23:chipyard.TestHarness.RocketConfig.fir@101385.4]
  wire [20:0] _T_1041; // @[Scheduler.scala 230:77:chipyard.TestHarness.RocketConfig.fir@101388.4]
  wire  _T_1044; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101391.4]
  wire [15:0] _GEN_148; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101392.4]
  wire [15:0] _T_1045; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101392.4]
  wire  _T_1048; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101395.4]
  wire [7:0] _T_1049; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101396.4]
  wire  _T_1052; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101399.4]
  wire [3:0] _T_1053; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101400.4]
  wire  _T_1056; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101403.4]
  wire [1:0] _T_1057; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101404.4]
  wire [3:0] _T_1061; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101408.4]
  wire  mshr_uses_directory_for_lb; // @[Scheduler.scala 237:45:chipyard.TestHarness.RocketConfig.fir@101415.4]
  wire [11:0] _T_1063; // @[Scheduler.scala 238:63:chipyard.TestHarness.RocketConfig.fir@101416.4]
  wire  _T_1064; // @[Scheduler.scala 238:56:chipyard.TestHarness.RocketConfig.fir@101417.4]
  wire  mshr_uses_directory; // @[Scheduler.scala 238:41:chipyard.TestHarness.RocketConfig.fir@101418.4]
  wire  alloc_uses_directory; // @[Scheduler.scala 251:44:chipyard.TestHarness.RocketConfig.fir@101448.4]
  wire  _T_1093; // @[Scheduler.scala 259:55:chipyard.TestHarness.RocketConfig.fir@101456.4]
  wire  _T_1098; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101463.4]
  wire [3:0] _GEN_149; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101464.4]
  wire [3:0] _T_1099; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101464.4]
  wire  _T_1102; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101467.4]
  wire [1:0] _T_1103; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101468.4]
  wire [2:0] _T_1106; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101471.4]
  wire [20:0] _T_1124; // @[Scheduler.scala 265:30:chipyard.TestHarness.RocketConfig.fir@101489.4]
  wire  _T_1127; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101492.4]
  wire [15:0] _GEN_151; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101493.4]
  wire [15:0] _T_1128; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101493.4]
  wire  _T_1131; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101496.4]
  wire [7:0] _T_1132; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101497.4]
  wire  _T_1135; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101500.4]
  wire [3:0] _T_1136; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101501.4]
  wire  _T_1139; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101504.4]
  wire [1:0] _T_1140; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101505.4]
  wire [4:0] _T_1145; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101510.4]
  wire [2:0] _T_1146; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101511.4]
  wire [4:0] _T_1148; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101513.4]
  wire [3:0] _T_1149; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101514.4]
  wire [4:0] _GEN_152; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101515.4]
  wire [7:0] _T_1153; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@101520.4]
  wire [6:0] _T_1155; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@101522.4]
  wire [8:0] _T_1156; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@101523.4]
  wire [6:0] _T_1158; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@101525.4]
  wire [10:0] _T_1159; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@101526.4]
  wire [6:0] _T_1161; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@101528.4]
  wire [7:0] _T_1163; // @[Scheduler.scala 267:47:chipyard.TestHarness.RocketConfig.fir@101530.4]
  wire [7:0] _T_1164; // @[Scheduler.scala 267:23:chipyard.TestHarness.RocketConfig.fir@101531.4]
  wire [7:0] _GEN_153; // @[Scheduler.scala 267:53:chipyard.TestHarness.RocketConfig.fir@101533.4]
  wire [7:0] _T_1166; // @[Scheduler.scala 267:53:chipyard.TestHarness.RocketConfig.fir@101533.4]
  wire [7:0] _GEN_154; // @[Scheduler.scala 267:69:chipyard.TestHarness.RocketConfig.fir@101534.4]
  wire [7:0] mshr_insertOH; // @[Scheduler.scala 267:69:chipyard.TestHarness.RocketConfig.fir@101534.4]
  wire  _T_1175; // @[Scheduler.scala 269:25:chipyard.TestHarness.RocketConfig.fir@101543.4]
  wire  _T_1176; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101544.4]
  wire  _T_1178; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101546.4]
  wire  _T_1180; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101553.4]
  wire  _T_1182; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101555.4]
  wire  _T_1184; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101562.4]
  wire  _T_1186; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101564.4]
  wire  _T_1188; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101571.4]
  wire  _T_1190; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101573.4]
  wire  _T_1192; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101580.4]
  wire  _T_1194; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101582.4]
  wire  _T_1196; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101589.4]
  wire  _T_1198; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101591.4]
  wire  _T_1200; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101598.4]
  wire  _T_1202; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101600.4]
  wire  _GEN_85; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  wire  _GEN_88; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  wire  _GEN_89; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  wire [2:0] _GEN_90; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  wire [2:0] _GEN_91; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  wire [2:0] _GEN_92; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  wire [2:0] _GEN_93; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  wire [11:0] _GEN_94; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  wire [5:0] _GEN_95; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  wire [5:0] _GEN_96; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  wire [9:0] _GEN_97; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  wire  _GEN_98; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  wire  _T_1212; // @[Scheduler.scala 280:12:chipyard.TestHarness.RocketConfig.fir@101619.6]
  wire  _T_1213; // @[Scheduler.scala 280:12:chipyard.TestHarness.RocketConfig.fir@101620.6]
  wire  _T_1216; // @[Scheduler.scala 284:32:chipyard.TestHarness.RocketConfig.fir@101629.4]
  wire  _T_1218; // @[Scheduler.scala 284:59:chipyard.TestHarness.RocketConfig.fir@101631.4]
  reg [7:0] directoryFanout; // @[Scheduler.scala 296:46:chipyard.TestHarness.RocketConfig.fir@101659.4]
  reg [31:0] _RAND_1;
  wire  _T_1237; // @[Scheduler.scala 304:63:chipyard.TestHarness.RocketConfig.fir@101682.4]
  wire  _T_1238; // @[Scheduler.scala 304:33:chipyard.TestHarness.RocketConfig.fir@101683.4]
  wire  _T_1239; // @[Scheduler.scala 306:74:chipyard.TestHarness.RocketConfig.fir@101684.4]
  wire  _T_1240; // @[Scheduler.scala 306:50:chipyard.TestHarness.RocketConfig.fir@101685.4]
  wire  _T_1241; // @[Scheduler.scala 306:74:chipyard.TestHarness.RocketConfig.fir@101686.4]
  wire  _T_1242; // @[Scheduler.scala 306:50:chipyard.TestHarness.RocketConfig.fir@101687.4]
  wire  _T_1243; // @[Scheduler.scala 306:74:chipyard.TestHarness.RocketConfig.fir@101688.4]
  wire  _T_1244; // @[Scheduler.scala 306:50:chipyard.TestHarness.RocketConfig.fir@101689.4]
  wire  _T_1245; // @[Scheduler.scala 306:74:chipyard.TestHarness.RocketConfig.fir@101690.4]
  wire  _T_1246; // @[Scheduler.scala 306:50:chipyard.TestHarness.RocketConfig.fir@101691.4]
  wire  _T_1247; // @[Scheduler.scala 306:74:chipyard.TestHarness.RocketConfig.fir@101692.4]
  wire  _T_1248; // @[Scheduler.scala 306:50:chipyard.TestHarness.RocketConfig.fir@101693.4]
  wire [2:0] _T_1249; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101694.4]
  wire [2:0] _T_1250; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101695.4]
  wire [2:0] _T_1251; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101696.4]
  wire [2:0] _T_1252; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101697.4]
  wire [2:0] _T_1253; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101698.4]
  wire [2:0] _T_1254; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101699.4]
  wire [2:0] _T_1255; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101700.4]
  wire [2:0] _T_1256; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101701.4]
  wire [2:0] _T_1257; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101702.4]
  wire [2:0] _T_1260_0; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101709.4]
  wire [2:0] _T_1260_1; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101710.4]
  wire [2:0] _GEN_128; // @[Scheduler.scala 308:16:chipyard.TestHarness.RocketConfig.fir@101716.4]
  wire [2:0] _T_1260_2; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101711.4]
  wire [2:0] _GEN_129; // @[Scheduler.scala 308:16:chipyard.TestHarness.RocketConfig.fir@101716.4]
  wire [2:0] _T_1260_3; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101712.4]
  wire [2:0] _GEN_130; // @[Scheduler.scala 308:16:chipyard.TestHarness.RocketConfig.fir@101716.4]
  wire [2:0] _T_1260_4; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101713.4]
  wire [2:0] _GEN_131; // @[Scheduler.scala 308:16:chipyard.TestHarness.RocketConfig.fir@101716.4]
  wire [2:0] _T_1260_5; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101714.4]
  wire [2:0] _GEN_132; // @[Scheduler.scala 308:16:chipyard.TestHarness.RocketConfig.fir@101716.4]
  wire [2:0] _T_1260_6; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101715.4]
  wire [9:0] _T_1261_0; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101719.4]
  wire [9:0] _T_1261_1; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101720.4]
  wire [9:0] _GEN_135; // @[Scheduler.scala 309:16:chipyard.TestHarness.RocketConfig.fir@101726.4]
  wire [9:0] _T_1261_2; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101721.4]
  wire [9:0] _GEN_136; // @[Scheduler.scala 309:16:chipyard.TestHarness.RocketConfig.fir@101726.4]
  wire [9:0] _T_1261_3; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101722.4]
  wire [9:0] _GEN_137; // @[Scheduler.scala 309:16:chipyard.TestHarness.RocketConfig.fir@101726.4]
  wire [9:0] _T_1261_4; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101723.4]
  wire [9:0] _GEN_138; // @[Scheduler.scala 309:16:chipyard.TestHarness.RocketConfig.fir@101726.4]
  wire [9:0] _T_1261_5; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101724.4]
  wire [9:0] _GEN_139; // @[Scheduler.scala 309:16:chipyard.TestHarness.RocketConfig.fir@101726.4]
  wire [9:0] _T_1261_6; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101725.4]
  SourceA sourceA ( // @[Scheduler.scala 38:23:chipyard.TestHarness.RocketConfig.fir@100029.4]
    .clock(sourceA_clock),
    .reset(sourceA_reset),
    .io_req_ready(sourceA_io_req_ready),
    .io_req_valid(sourceA_io_req_valid),
    .io_req_bits_tag(sourceA_io_req_bits_tag),
    .io_req_bits_set(sourceA_io_req_bits_set),
    .io_req_bits_param(sourceA_io_req_bits_param),
    .io_req_bits_source(sourceA_io_req_bits_source),
    .io_req_bits_block(sourceA_io_req_bits_block),
    .io_a_ready(sourceA_io_a_ready),
    .io_a_valid(sourceA_io_a_valid),
    .io_a_bits_opcode(sourceA_io_a_bits_opcode),
    .io_a_bits_param(sourceA_io_a_bits_param),
    .io_a_bits_size(sourceA_io_a_bits_size),
    .io_a_bits_source(sourceA_io_a_bits_source),
    .io_a_bits_address(sourceA_io_a_bits_address),
    .io_a_bits_mask(sourceA_io_a_bits_mask),
    .io_a_bits_data(sourceA_io_a_bits_data),
    .io_a_bits_corrupt(sourceA_io_a_bits_corrupt)
  );
  SourceB sourceB ( // @[Scheduler.scala 39:23:chipyard.TestHarness.RocketConfig.fir@100033.4]
    .clock(sourceB_clock),
    .reset(sourceB_reset),
    .io_req_ready(sourceB_io_req_ready),
    .io_req_valid(sourceB_io_req_valid),
    .io_req_bits_param(sourceB_io_req_bits_param),
    .io_req_bits_tag(sourceB_io_req_bits_tag),
    .io_req_bits_set(sourceB_io_req_bits_set),
    .io_req_bits_clients(sourceB_io_req_bits_clients),
    .io_b_ready(sourceB_io_b_ready),
    .io_b_valid(sourceB_io_b_valid),
    .io_b_bits_param(sourceB_io_b_bits_param),
    .io_b_bits_address(sourceB_io_b_bits_address)
  );
  SourceC sourceC ( // @[Scheduler.scala 40:23:chipyard.TestHarness.RocketConfig.fir@100037.4]
    .clock(sourceC_clock),
    .reset(sourceC_reset),
    .io_req_ready(sourceC_io_req_ready),
    .io_req_valid(sourceC_io_req_valid),
    .io_req_bits_opcode(sourceC_io_req_bits_opcode),
    .io_req_bits_param(sourceC_io_req_bits_param),
    .io_req_bits_source(sourceC_io_req_bits_source),
    .io_req_bits_tag(sourceC_io_req_bits_tag),
    .io_req_bits_set(sourceC_io_req_bits_set),
    .io_req_bits_way(sourceC_io_req_bits_way),
    .io_req_bits_dirty(sourceC_io_req_bits_dirty),
    .io_c_ready(sourceC_io_c_ready),
    .io_c_valid(sourceC_io_c_valid),
    .io_c_bits_opcode(sourceC_io_c_bits_opcode),
    .io_c_bits_param(sourceC_io_c_bits_param),
    .io_c_bits_size(sourceC_io_c_bits_size),
    .io_c_bits_source(sourceC_io_c_bits_source),
    .io_c_bits_address(sourceC_io_c_bits_address),
    .io_c_bits_data(sourceC_io_c_bits_data),
    .io_c_bits_corrupt(sourceC_io_c_bits_corrupt),
    .io_bs_adr_ready(sourceC_io_bs_adr_ready),
    .io_bs_adr_valid(sourceC_io_bs_adr_valid),
    .io_bs_adr_bits_way(sourceC_io_bs_adr_bits_way),
    .io_bs_adr_bits_set(sourceC_io_bs_adr_bits_set),
    .io_bs_adr_bits_beat(sourceC_io_bs_adr_bits_beat),
    .io_bs_dat_data(sourceC_io_bs_dat_data),
    .io_evict_req_set(sourceC_io_evict_req_set),
    .io_evict_req_way(sourceC_io_evict_req_way),
    .io_evict_safe(sourceC_io_evict_safe)
  );
  SourceD sourceD ( // @[Scheduler.scala 41:23:chipyard.TestHarness.RocketConfig.fir@100041.4]
    .clock(sourceD_clock),
    .reset(sourceD_reset),
    .io_req_ready(sourceD_io_req_ready),
    .io_req_valid(sourceD_io_req_valid),
    .io_req_bits_prio_0(sourceD_io_req_bits_prio_0),
    .io_req_bits_prio_2(sourceD_io_req_bits_prio_2),
    .io_req_bits_opcode(sourceD_io_req_bits_opcode),
    .io_req_bits_param(sourceD_io_req_bits_param),
    .io_req_bits_size(sourceD_io_req_bits_size),
    .io_req_bits_source(sourceD_io_req_bits_source),
    .io_req_bits_offset(sourceD_io_req_bits_offset),
    .io_req_bits_put(sourceD_io_req_bits_put),
    .io_req_bits_set(sourceD_io_req_bits_set),
    .io_req_bits_sink(sourceD_io_req_bits_sink),
    .io_req_bits_way(sourceD_io_req_bits_way),
    .io_req_bits_bad(sourceD_io_req_bits_bad),
    .io_d_ready(sourceD_io_d_ready),
    .io_d_valid(sourceD_io_d_valid),
    .io_d_bits_opcode(sourceD_io_d_bits_opcode),
    .io_d_bits_param(sourceD_io_d_bits_param),
    .io_d_bits_size(sourceD_io_d_bits_size),
    .io_d_bits_source(sourceD_io_d_bits_source),
    .io_d_bits_sink(sourceD_io_d_bits_sink),
    .io_d_bits_denied(sourceD_io_d_bits_denied),
    .io_d_bits_data(sourceD_io_d_bits_data),
    .io_d_bits_corrupt(sourceD_io_d_bits_corrupt),
    .io_pb_pop_ready(sourceD_io_pb_pop_ready),
    .io_pb_pop_valid(sourceD_io_pb_pop_valid),
    .io_pb_pop_bits_index(sourceD_io_pb_pop_bits_index),
    .io_pb_pop_bits_last(sourceD_io_pb_pop_bits_last),
    .io_pb_beat_data(sourceD_io_pb_beat_data),
    .io_pb_beat_mask(sourceD_io_pb_beat_mask),
    .io_pb_beat_corrupt(sourceD_io_pb_beat_corrupt),
    .io_rel_pop_ready(sourceD_io_rel_pop_ready),
    .io_rel_pop_valid(sourceD_io_rel_pop_valid),
    .io_rel_pop_bits_index(sourceD_io_rel_pop_bits_index),
    .io_rel_pop_bits_last(sourceD_io_rel_pop_bits_last),
    .io_rel_beat_data(sourceD_io_rel_beat_data),
    .io_rel_beat_corrupt(sourceD_io_rel_beat_corrupt),
    .io_bs_radr_ready(sourceD_io_bs_radr_ready),
    .io_bs_radr_valid(sourceD_io_bs_radr_valid),
    .io_bs_radr_bits_way(sourceD_io_bs_radr_bits_way),
    .io_bs_radr_bits_set(sourceD_io_bs_radr_bits_set),
    .io_bs_radr_bits_beat(sourceD_io_bs_radr_bits_beat),
    .io_bs_radr_bits_mask(sourceD_io_bs_radr_bits_mask),
    .io_bs_rdat_data(sourceD_io_bs_rdat_data),
    .io_bs_wadr_ready(sourceD_io_bs_wadr_ready),
    .io_bs_wadr_valid(sourceD_io_bs_wadr_valid),
    .io_bs_wadr_bits_way(sourceD_io_bs_wadr_bits_way),
    .io_bs_wadr_bits_set(sourceD_io_bs_wadr_bits_set),
    .io_bs_wadr_bits_beat(sourceD_io_bs_wadr_bits_beat),
    .io_bs_wadr_bits_mask(sourceD_io_bs_wadr_bits_mask),
    .io_bs_wdat_data(sourceD_io_bs_wdat_data),
    .io_evict_req_set(sourceD_io_evict_req_set),
    .io_evict_req_way(sourceD_io_evict_req_way),
    .io_evict_safe(sourceD_io_evict_safe),
    .io_grant_req_set(sourceD_io_grant_req_set),
    .io_grant_req_way(sourceD_io_grant_req_way),
    .io_grant_safe(sourceD_io_grant_safe)
  );
  SourceE sourceE ( // @[Scheduler.scala 42:23:chipyard.TestHarness.RocketConfig.fir@100045.4]
    .clock(sourceE_clock),
    .reset(sourceE_reset),
    .io_req_ready(sourceE_io_req_ready),
    .io_req_valid(sourceE_io_req_valid),
    .io_req_bits_sink(sourceE_io_req_bits_sink),
    .io_e_valid(sourceE_io_e_valid),
    .io_e_bits_sink(sourceE_io_e_bits_sink)
  );
  SourceX sourceX ( // @[Scheduler.scala 43:23:chipyard.TestHarness.RocketConfig.fir@100049.4]
    .clock(sourceX_clock),
    .reset(sourceX_reset),
    .io_req_ready(sourceX_io_req_ready),
    .io_req_valid(sourceX_io_req_valid),
    .io_x_ready(sourceX_io_x_ready),
    .io_x_valid(sourceX_io_x_valid)
  );
  SinkA sinkA ( // @[Scheduler.scala 52:21:chipyard.TestHarness.RocketConfig.fir@100059.4]
    .clock(sinkA_clock),
    .reset(sinkA_reset),
    .io_req_ready(sinkA_io_req_ready),
    .io_req_valid(sinkA_io_req_valid),
    .io_req_bits_opcode(sinkA_io_req_bits_opcode),
    .io_req_bits_param(sinkA_io_req_bits_param),
    .io_req_bits_size(sinkA_io_req_bits_size),
    .io_req_bits_source(sinkA_io_req_bits_source),
    .io_req_bits_tag(sinkA_io_req_bits_tag),
    .io_req_bits_offset(sinkA_io_req_bits_offset),
    .io_req_bits_put(sinkA_io_req_bits_put),
    .io_req_bits_set(sinkA_io_req_bits_set),
    .io_a_ready(sinkA_io_a_ready),
    .io_a_valid(sinkA_io_a_valid),
    .io_a_bits_opcode(sinkA_io_a_bits_opcode),
    .io_a_bits_param(sinkA_io_a_bits_param),
    .io_a_bits_size(sinkA_io_a_bits_size),
    .io_a_bits_source(sinkA_io_a_bits_source),
    .io_a_bits_address(sinkA_io_a_bits_address),
    .io_a_bits_mask(sinkA_io_a_bits_mask),
    .io_a_bits_data(sinkA_io_a_bits_data),
    .io_a_bits_corrupt(sinkA_io_a_bits_corrupt),
    .io_pb_pop_ready(sinkA_io_pb_pop_ready),
    .io_pb_pop_valid(sinkA_io_pb_pop_valid),
    .io_pb_pop_bits_index(sinkA_io_pb_pop_bits_index),
    .io_pb_pop_bits_last(sinkA_io_pb_pop_bits_last),
    .io_pb_beat_data(sinkA_io_pb_beat_data),
    .io_pb_beat_mask(sinkA_io_pb_beat_mask),
    .io_pb_beat_corrupt(sinkA_io_pb_beat_corrupt)
  );
  SinkC sinkC ( // @[Scheduler.scala 53:21:chipyard.TestHarness.RocketConfig.fir@100063.4]
    .clock(sinkC_clock),
    .reset(sinkC_reset),
    .io_req_ready(sinkC_io_req_ready),
    .io_req_valid(sinkC_io_req_valid),
    .io_req_bits_opcode(sinkC_io_req_bits_opcode),
    .io_req_bits_param(sinkC_io_req_bits_param),
    .io_req_bits_size(sinkC_io_req_bits_size),
    .io_req_bits_source(sinkC_io_req_bits_source),
    .io_req_bits_tag(sinkC_io_req_bits_tag),
    .io_req_bits_offset(sinkC_io_req_bits_offset),
    .io_req_bits_put(sinkC_io_req_bits_put),
    .io_req_bits_set(sinkC_io_req_bits_set),
    .io_resp_valid(sinkC_io_resp_valid),
    .io_resp_bits_last(sinkC_io_resp_bits_last),
    .io_resp_bits_set(sinkC_io_resp_bits_set),
    .io_resp_bits_tag(sinkC_io_resp_bits_tag),
    .io_resp_bits_source(sinkC_io_resp_bits_source),
    .io_resp_bits_param(sinkC_io_resp_bits_param),
    .io_resp_bits_data(sinkC_io_resp_bits_data),
    .io_c_ready(sinkC_io_c_ready),
    .io_c_valid(sinkC_io_c_valid),
    .io_c_bits_opcode(sinkC_io_c_bits_opcode),
    .io_c_bits_param(sinkC_io_c_bits_param),
    .io_c_bits_size(sinkC_io_c_bits_size),
    .io_c_bits_source(sinkC_io_c_bits_source),
    .io_c_bits_address(sinkC_io_c_bits_address),
    .io_c_bits_data(sinkC_io_c_bits_data),
    .io_c_bits_corrupt(sinkC_io_c_bits_corrupt),
    .io_set(sinkC_io_set),
    .io_way(sinkC_io_way),
    .io_bs_adr_ready(sinkC_io_bs_adr_ready),
    .io_bs_adr_valid(sinkC_io_bs_adr_valid),
    .io_bs_adr_bits_noop(sinkC_io_bs_adr_bits_noop),
    .io_bs_adr_bits_way(sinkC_io_bs_adr_bits_way),
    .io_bs_adr_bits_set(sinkC_io_bs_adr_bits_set),
    .io_bs_adr_bits_beat(sinkC_io_bs_adr_bits_beat),
    .io_bs_adr_bits_mask(sinkC_io_bs_adr_bits_mask),
    .io_bs_dat_data(sinkC_io_bs_dat_data),
    .io_rel_pop_ready(sinkC_io_rel_pop_ready),
    .io_rel_pop_valid(sinkC_io_rel_pop_valid),
    .io_rel_pop_bits_index(sinkC_io_rel_pop_bits_index),
    .io_rel_pop_bits_last(sinkC_io_rel_pop_bits_last),
    .io_rel_beat_data(sinkC_io_rel_beat_data),
    .io_rel_beat_corrupt(sinkC_io_rel_beat_corrupt)
  );
  SinkD sinkD ( // @[Scheduler.scala 54:21:chipyard.TestHarness.RocketConfig.fir@100067.4]
    .clock(sinkD_clock),
    .reset(sinkD_reset),
    .io_resp_valid(sinkD_io_resp_valid),
    .io_resp_bits_last(sinkD_io_resp_bits_last),
    .io_resp_bits_opcode(sinkD_io_resp_bits_opcode),
    .io_resp_bits_param(sinkD_io_resp_bits_param),
    .io_resp_bits_source(sinkD_io_resp_bits_source),
    .io_resp_bits_sink(sinkD_io_resp_bits_sink),
    .io_resp_bits_denied(sinkD_io_resp_bits_denied),
    .io_d_ready(sinkD_io_d_ready),
    .io_d_valid(sinkD_io_d_valid),
    .io_d_bits_opcode(sinkD_io_d_bits_opcode),
    .io_d_bits_param(sinkD_io_d_bits_param),
    .io_d_bits_size(sinkD_io_d_bits_size),
    .io_d_bits_source(sinkD_io_d_bits_source),
    .io_d_bits_sink(sinkD_io_d_bits_sink),
    .io_d_bits_denied(sinkD_io_d_bits_denied),
    .io_d_bits_data(sinkD_io_d_bits_data),
    .io_d_bits_corrupt(sinkD_io_d_bits_corrupt),
    .io_source(sinkD_io_source),
    .io_way(sinkD_io_way),
    .io_set(sinkD_io_set),
    .io_bs_adr_ready(sinkD_io_bs_adr_ready),
    .io_bs_adr_valid(sinkD_io_bs_adr_valid),
    .io_bs_adr_bits_noop(sinkD_io_bs_adr_bits_noop),
    .io_bs_adr_bits_way(sinkD_io_bs_adr_bits_way),
    .io_bs_adr_bits_set(sinkD_io_bs_adr_bits_set),
    .io_bs_adr_bits_beat(sinkD_io_bs_adr_bits_beat),
    .io_bs_dat_data(sinkD_io_bs_dat_data),
    .io_grant_req_set(sinkD_io_grant_req_set),
    .io_grant_req_way(sinkD_io_grant_req_way),
    .io_grant_safe(sinkD_io_grant_safe)
  );
  SinkE sinkE ( // @[Scheduler.scala 55:21:chipyard.TestHarness.RocketConfig.fir@100071.4]
    .io_resp_valid(sinkE_io_resp_valid),
    .io_resp_bits_sink(sinkE_io_resp_bits_sink),
    .io_e_valid(sinkE_io_e_valid),
    .io_e_bits_sink(sinkE_io_e_bits_sink)
  );
  SinkX sinkX ( // @[Scheduler.scala 56:21:chipyard.TestHarness.RocketConfig.fir@100075.4]
    .clock(sinkX_clock),
    .reset(sinkX_reset),
    .io_req_ready(sinkX_io_req_ready),
    .io_req_valid(sinkX_io_req_valid),
    .io_req_bits_tag(sinkX_io_req_bits_tag),
    .io_req_bits_set(sinkX_io_req_bits_set),
    .io_x_ready(sinkX_io_x_ready),
    .io_x_valid(sinkX_io_x_valid),
    .io_x_bits_address(sinkX_io_x_bits_address)
  );
  Directory directory ( // @[Scheduler.scala 66:25:chipyard.TestHarness.RocketConfig.fir@100085.4]
    .clock(directory_clock),
    .reset(directory_reset),
    .io_write_ready(directory_io_write_ready),
    .io_write_valid(directory_io_write_valid),
    .io_write_bits_set(directory_io_write_bits_set),
    .io_write_bits_way(directory_io_write_bits_way),
    .io_write_bits_data_dirty(directory_io_write_bits_data_dirty),
    .io_write_bits_data_state(directory_io_write_bits_data_state),
    .io_write_bits_data_clients(directory_io_write_bits_data_clients),
    .io_write_bits_data_tag(directory_io_write_bits_data_tag),
    .io_read_valid(directory_io_read_valid),
    .io_read_bits_set(directory_io_read_bits_set),
    .io_read_bits_tag(directory_io_read_bits_tag),
    .io_result_bits_dirty(directory_io_result_bits_dirty),
    .io_result_bits_state(directory_io_result_bits_state),
    .io_result_bits_clients(directory_io_result_bits_clients),
    .io_result_bits_tag(directory_io_result_bits_tag),
    .io_result_bits_hit(directory_io_result_bits_hit),
    .io_result_bits_way(directory_io_result_bits_way),
    .io_ready(directory_io_ready)
  );
  BankedStore bankedStore ( // @[Scheduler.scala 67:27:chipyard.TestHarness.RocketConfig.fir@100089.4]
    .clock(bankedStore_clock),
    .io_sinkC_adr_ready(bankedStore_io_sinkC_adr_ready),
    .io_sinkC_adr_valid(bankedStore_io_sinkC_adr_valid),
    .io_sinkC_adr_bits_noop(bankedStore_io_sinkC_adr_bits_noop),
    .io_sinkC_adr_bits_way(bankedStore_io_sinkC_adr_bits_way),
    .io_sinkC_adr_bits_set(bankedStore_io_sinkC_adr_bits_set),
    .io_sinkC_adr_bits_beat(bankedStore_io_sinkC_adr_bits_beat),
    .io_sinkC_adr_bits_mask(bankedStore_io_sinkC_adr_bits_mask),
    .io_sinkC_dat_data(bankedStore_io_sinkC_dat_data),
    .io_sinkD_adr_ready(bankedStore_io_sinkD_adr_ready),
    .io_sinkD_adr_valid(bankedStore_io_sinkD_adr_valid),
    .io_sinkD_adr_bits_noop(bankedStore_io_sinkD_adr_bits_noop),
    .io_sinkD_adr_bits_way(bankedStore_io_sinkD_adr_bits_way),
    .io_sinkD_adr_bits_set(bankedStore_io_sinkD_adr_bits_set),
    .io_sinkD_adr_bits_beat(bankedStore_io_sinkD_adr_bits_beat),
    .io_sinkD_dat_data(bankedStore_io_sinkD_dat_data),
    .io_sourceC_adr_ready(bankedStore_io_sourceC_adr_ready),
    .io_sourceC_adr_valid(bankedStore_io_sourceC_adr_valid),
    .io_sourceC_adr_bits_way(bankedStore_io_sourceC_adr_bits_way),
    .io_sourceC_adr_bits_set(bankedStore_io_sourceC_adr_bits_set),
    .io_sourceC_adr_bits_beat(bankedStore_io_sourceC_adr_bits_beat),
    .io_sourceC_dat_data(bankedStore_io_sourceC_dat_data),
    .io_sourceD_radr_ready(bankedStore_io_sourceD_radr_ready),
    .io_sourceD_radr_valid(bankedStore_io_sourceD_radr_valid),
    .io_sourceD_radr_bits_way(bankedStore_io_sourceD_radr_bits_way),
    .io_sourceD_radr_bits_set(bankedStore_io_sourceD_radr_bits_set),
    .io_sourceD_radr_bits_beat(bankedStore_io_sourceD_radr_bits_beat),
    .io_sourceD_radr_bits_mask(bankedStore_io_sourceD_radr_bits_mask),
    .io_sourceD_rdat_data(bankedStore_io_sourceD_rdat_data),
    .io_sourceD_wadr_ready(bankedStore_io_sourceD_wadr_ready),
    .io_sourceD_wadr_valid(bankedStore_io_sourceD_wadr_valid),
    .io_sourceD_wadr_bits_way(bankedStore_io_sourceD_wadr_bits_way),
    .io_sourceD_wadr_bits_set(bankedStore_io_sourceD_wadr_bits_set),
    .io_sourceD_wadr_bits_beat(bankedStore_io_sourceD_wadr_bits_beat),
    .io_sourceD_wadr_bits_mask(bankedStore_io_sourceD_wadr_bits_mask),
    .io_sourceD_wdat_data(bankedStore_io_sourceD_wdat_data)
  );
  ListBuffer_2 requests ( // @[Scheduler.scala 68:24:chipyard.TestHarness.RocketConfig.fir@100093.4]
    .clock(requests_clock),
    .reset(requests_reset),
    .io_push_ready(requests_io_push_ready),
    .io_push_valid(requests_io_push_valid),
    .io_push_bits_index(requests_io_push_bits_index),
    .io_push_bits_data_prio_0(requests_io_push_bits_data_prio_0),
    .io_push_bits_data_prio_2(requests_io_push_bits_data_prio_2),
    .io_push_bits_data_control(requests_io_push_bits_data_control),
    .io_push_bits_data_opcode(requests_io_push_bits_data_opcode),
    .io_push_bits_data_param(requests_io_push_bits_data_param),
    .io_push_bits_data_size(requests_io_push_bits_data_size),
    .io_push_bits_data_source(requests_io_push_bits_data_source),
    .io_push_bits_data_tag(requests_io_push_bits_data_tag),
    .io_push_bits_data_offset(requests_io_push_bits_data_offset),
    .io_push_bits_data_put(requests_io_push_bits_data_put),
    .io_valid(requests_io_valid),
    .io_pop_valid(requests_io_pop_valid),
    .io_pop_bits(requests_io_pop_bits),
    .io_data_prio_0(requests_io_data_prio_0),
    .io_data_prio_1(requests_io_data_prio_1),
    .io_data_prio_2(requests_io_data_prio_2),
    .io_data_control(requests_io_data_control),
    .io_data_opcode(requests_io_data_opcode),
    .io_data_param(requests_io_data_param),
    .io_data_size(requests_io_data_size),
    .io_data_source(requests_io_data_source),
    .io_data_tag(requests_io_data_tag),
    .io_data_offset(requests_io_data_offset),
    .io_data_put(requests_io_data_put)
  );
  MSHR abc_mshrs_0 ( // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100097.4]
    .clock(abc_mshrs_0_clock),
    .reset(abc_mshrs_0_reset),
    .io_allocate_valid(abc_mshrs_0_io_allocate_valid),
    .io_allocate_bits_prio_0(abc_mshrs_0_io_allocate_bits_prio_0),
    .io_allocate_bits_prio_1(abc_mshrs_0_io_allocate_bits_prio_1),
    .io_allocate_bits_prio_2(abc_mshrs_0_io_allocate_bits_prio_2),
    .io_allocate_bits_control(abc_mshrs_0_io_allocate_bits_control),
    .io_allocate_bits_opcode(abc_mshrs_0_io_allocate_bits_opcode),
    .io_allocate_bits_param(abc_mshrs_0_io_allocate_bits_param),
    .io_allocate_bits_size(abc_mshrs_0_io_allocate_bits_size),
    .io_allocate_bits_source(abc_mshrs_0_io_allocate_bits_source),
    .io_allocate_bits_tag(abc_mshrs_0_io_allocate_bits_tag),
    .io_allocate_bits_offset(abc_mshrs_0_io_allocate_bits_offset),
    .io_allocate_bits_put(abc_mshrs_0_io_allocate_bits_put),
    .io_allocate_bits_set(abc_mshrs_0_io_allocate_bits_set),
    .io_allocate_bits_repeat(abc_mshrs_0_io_allocate_bits_repeat),
    .io_directory_valid(abc_mshrs_0_io_directory_valid),
    .io_directory_bits_dirty(abc_mshrs_0_io_directory_bits_dirty),
    .io_directory_bits_state(abc_mshrs_0_io_directory_bits_state),
    .io_directory_bits_clients(abc_mshrs_0_io_directory_bits_clients),
    .io_directory_bits_tag(abc_mshrs_0_io_directory_bits_tag),
    .io_directory_bits_hit(abc_mshrs_0_io_directory_bits_hit),
    .io_directory_bits_way(abc_mshrs_0_io_directory_bits_way),
    .io_status_valid(abc_mshrs_0_io_status_valid),
    .io_status_bits_set(abc_mshrs_0_io_status_bits_set),
    .io_status_bits_tag(abc_mshrs_0_io_status_bits_tag),
    .io_status_bits_way(abc_mshrs_0_io_status_bits_way),
    .io_status_bits_blockB(abc_mshrs_0_io_status_bits_blockB),
    .io_status_bits_nestB(abc_mshrs_0_io_status_bits_nestB),
    .io_status_bits_blockC(abc_mshrs_0_io_status_bits_blockC),
    .io_status_bits_nestC(abc_mshrs_0_io_status_bits_nestC),
    .io_schedule_ready(abc_mshrs_0_io_schedule_ready),
    .io_schedule_valid(abc_mshrs_0_io_schedule_valid),
    .io_schedule_bits_a_valid(abc_mshrs_0_io_schedule_bits_a_valid),
    .io_schedule_bits_a_bits_tag(abc_mshrs_0_io_schedule_bits_a_bits_tag),
    .io_schedule_bits_a_bits_set(abc_mshrs_0_io_schedule_bits_a_bits_set),
    .io_schedule_bits_a_bits_param(abc_mshrs_0_io_schedule_bits_a_bits_param),
    .io_schedule_bits_a_bits_block(abc_mshrs_0_io_schedule_bits_a_bits_block),
    .io_schedule_bits_b_valid(abc_mshrs_0_io_schedule_bits_b_valid),
    .io_schedule_bits_b_bits_param(abc_mshrs_0_io_schedule_bits_b_bits_param),
    .io_schedule_bits_b_bits_tag(abc_mshrs_0_io_schedule_bits_b_bits_tag),
    .io_schedule_bits_b_bits_set(abc_mshrs_0_io_schedule_bits_b_bits_set),
    .io_schedule_bits_b_bits_clients(abc_mshrs_0_io_schedule_bits_b_bits_clients),
    .io_schedule_bits_c_valid(abc_mshrs_0_io_schedule_bits_c_valid),
    .io_schedule_bits_c_bits_opcode(abc_mshrs_0_io_schedule_bits_c_bits_opcode),
    .io_schedule_bits_c_bits_param(abc_mshrs_0_io_schedule_bits_c_bits_param),
    .io_schedule_bits_c_bits_tag(abc_mshrs_0_io_schedule_bits_c_bits_tag),
    .io_schedule_bits_c_bits_set(abc_mshrs_0_io_schedule_bits_c_bits_set),
    .io_schedule_bits_c_bits_way(abc_mshrs_0_io_schedule_bits_c_bits_way),
    .io_schedule_bits_c_bits_dirty(abc_mshrs_0_io_schedule_bits_c_bits_dirty),
    .io_schedule_bits_d_valid(abc_mshrs_0_io_schedule_bits_d_valid),
    .io_schedule_bits_d_bits_prio_0(abc_mshrs_0_io_schedule_bits_d_bits_prio_0),
    .io_schedule_bits_d_bits_prio_1(abc_mshrs_0_io_schedule_bits_d_bits_prio_1),
    .io_schedule_bits_d_bits_prio_2(abc_mshrs_0_io_schedule_bits_d_bits_prio_2),
    .io_schedule_bits_d_bits_control(abc_mshrs_0_io_schedule_bits_d_bits_control),
    .io_schedule_bits_d_bits_opcode(abc_mshrs_0_io_schedule_bits_d_bits_opcode),
    .io_schedule_bits_d_bits_param(abc_mshrs_0_io_schedule_bits_d_bits_param),
    .io_schedule_bits_d_bits_size(abc_mshrs_0_io_schedule_bits_d_bits_size),
    .io_schedule_bits_d_bits_source(abc_mshrs_0_io_schedule_bits_d_bits_source),
    .io_schedule_bits_d_bits_tag(abc_mshrs_0_io_schedule_bits_d_bits_tag),
    .io_schedule_bits_d_bits_offset(abc_mshrs_0_io_schedule_bits_d_bits_offset),
    .io_schedule_bits_d_bits_put(abc_mshrs_0_io_schedule_bits_d_bits_put),
    .io_schedule_bits_d_bits_set(abc_mshrs_0_io_schedule_bits_d_bits_set),
    .io_schedule_bits_d_bits_way(abc_mshrs_0_io_schedule_bits_d_bits_way),
    .io_schedule_bits_d_bits_bad(abc_mshrs_0_io_schedule_bits_d_bits_bad),
    .io_schedule_bits_e_valid(abc_mshrs_0_io_schedule_bits_e_valid),
    .io_schedule_bits_e_bits_sink(abc_mshrs_0_io_schedule_bits_e_bits_sink),
    .io_schedule_bits_x_valid(abc_mshrs_0_io_schedule_bits_x_valid),
    .io_schedule_bits_dir_valid(abc_mshrs_0_io_schedule_bits_dir_valid),
    .io_schedule_bits_dir_bits_set(abc_mshrs_0_io_schedule_bits_dir_bits_set),
    .io_schedule_bits_dir_bits_way(abc_mshrs_0_io_schedule_bits_dir_bits_way),
    .io_schedule_bits_dir_bits_data_dirty(abc_mshrs_0_io_schedule_bits_dir_bits_data_dirty),
    .io_schedule_bits_dir_bits_data_state(abc_mshrs_0_io_schedule_bits_dir_bits_data_state),
    .io_schedule_bits_dir_bits_data_clients(abc_mshrs_0_io_schedule_bits_dir_bits_data_clients),
    .io_schedule_bits_dir_bits_data_tag(abc_mshrs_0_io_schedule_bits_dir_bits_data_tag),
    .io_schedule_bits_reload(abc_mshrs_0_io_schedule_bits_reload),
    .io_sinkc_valid(abc_mshrs_0_io_sinkc_valid),
    .io_sinkc_bits_last(abc_mshrs_0_io_sinkc_bits_last),
    .io_sinkc_bits_tag(abc_mshrs_0_io_sinkc_bits_tag),
    .io_sinkc_bits_source(abc_mshrs_0_io_sinkc_bits_source),
    .io_sinkc_bits_param(abc_mshrs_0_io_sinkc_bits_param),
    .io_sinkc_bits_data(abc_mshrs_0_io_sinkc_bits_data),
    .io_sinkd_valid(abc_mshrs_0_io_sinkd_valid),
    .io_sinkd_bits_last(abc_mshrs_0_io_sinkd_bits_last),
    .io_sinkd_bits_opcode(abc_mshrs_0_io_sinkd_bits_opcode),
    .io_sinkd_bits_param(abc_mshrs_0_io_sinkd_bits_param),
    .io_sinkd_bits_sink(abc_mshrs_0_io_sinkd_bits_sink),
    .io_sinkd_bits_denied(abc_mshrs_0_io_sinkd_bits_denied),
    .io_sinke_valid(abc_mshrs_0_io_sinke_valid),
    .io_nestedwb_set(abc_mshrs_0_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshrs_0_io_nestedwb_tag),
    .io_nestedwb_b_toN(abc_mshrs_0_io_nestedwb_b_toN),
    .io_nestedwb_b_toB(abc_mshrs_0_io_nestedwb_b_toB),
    .io_nestedwb_b_clr_dirty(abc_mshrs_0_io_nestedwb_b_clr_dirty),
    .io_nestedwb_c_set_dirty(abc_mshrs_0_io_nestedwb_c_set_dirty)
  );
  MSHR abc_mshrs_1 ( // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100101.4]
    .clock(abc_mshrs_1_clock),
    .reset(abc_mshrs_1_reset),
    .io_allocate_valid(abc_mshrs_1_io_allocate_valid),
    .io_allocate_bits_prio_0(abc_mshrs_1_io_allocate_bits_prio_0),
    .io_allocate_bits_prio_1(abc_mshrs_1_io_allocate_bits_prio_1),
    .io_allocate_bits_prio_2(abc_mshrs_1_io_allocate_bits_prio_2),
    .io_allocate_bits_control(abc_mshrs_1_io_allocate_bits_control),
    .io_allocate_bits_opcode(abc_mshrs_1_io_allocate_bits_opcode),
    .io_allocate_bits_param(abc_mshrs_1_io_allocate_bits_param),
    .io_allocate_bits_size(abc_mshrs_1_io_allocate_bits_size),
    .io_allocate_bits_source(abc_mshrs_1_io_allocate_bits_source),
    .io_allocate_bits_tag(abc_mshrs_1_io_allocate_bits_tag),
    .io_allocate_bits_offset(abc_mshrs_1_io_allocate_bits_offset),
    .io_allocate_bits_put(abc_mshrs_1_io_allocate_bits_put),
    .io_allocate_bits_set(abc_mshrs_1_io_allocate_bits_set),
    .io_allocate_bits_repeat(abc_mshrs_1_io_allocate_bits_repeat),
    .io_directory_valid(abc_mshrs_1_io_directory_valid),
    .io_directory_bits_dirty(abc_mshrs_1_io_directory_bits_dirty),
    .io_directory_bits_state(abc_mshrs_1_io_directory_bits_state),
    .io_directory_bits_clients(abc_mshrs_1_io_directory_bits_clients),
    .io_directory_bits_tag(abc_mshrs_1_io_directory_bits_tag),
    .io_directory_bits_hit(abc_mshrs_1_io_directory_bits_hit),
    .io_directory_bits_way(abc_mshrs_1_io_directory_bits_way),
    .io_status_valid(abc_mshrs_1_io_status_valid),
    .io_status_bits_set(abc_mshrs_1_io_status_bits_set),
    .io_status_bits_tag(abc_mshrs_1_io_status_bits_tag),
    .io_status_bits_way(abc_mshrs_1_io_status_bits_way),
    .io_status_bits_blockB(abc_mshrs_1_io_status_bits_blockB),
    .io_status_bits_nestB(abc_mshrs_1_io_status_bits_nestB),
    .io_status_bits_blockC(abc_mshrs_1_io_status_bits_blockC),
    .io_status_bits_nestC(abc_mshrs_1_io_status_bits_nestC),
    .io_schedule_ready(abc_mshrs_1_io_schedule_ready),
    .io_schedule_valid(abc_mshrs_1_io_schedule_valid),
    .io_schedule_bits_a_valid(abc_mshrs_1_io_schedule_bits_a_valid),
    .io_schedule_bits_a_bits_tag(abc_mshrs_1_io_schedule_bits_a_bits_tag),
    .io_schedule_bits_a_bits_set(abc_mshrs_1_io_schedule_bits_a_bits_set),
    .io_schedule_bits_a_bits_param(abc_mshrs_1_io_schedule_bits_a_bits_param),
    .io_schedule_bits_a_bits_block(abc_mshrs_1_io_schedule_bits_a_bits_block),
    .io_schedule_bits_b_valid(abc_mshrs_1_io_schedule_bits_b_valid),
    .io_schedule_bits_b_bits_param(abc_mshrs_1_io_schedule_bits_b_bits_param),
    .io_schedule_bits_b_bits_tag(abc_mshrs_1_io_schedule_bits_b_bits_tag),
    .io_schedule_bits_b_bits_set(abc_mshrs_1_io_schedule_bits_b_bits_set),
    .io_schedule_bits_b_bits_clients(abc_mshrs_1_io_schedule_bits_b_bits_clients),
    .io_schedule_bits_c_valid(abc_mshrs_1_io_schedule_bits_c_valid),
    .io_schedule_bits_c_bits_opcode(abc_mshrs_1_io_schedule_bits_c_bits_opcode),
    .io_schedule_bits_c_bits_param(abc_mshrs_1_io_schedule_bits_c_bits_param),
    .io_schedule_bits_c_bits_tag(abc_mshrs_1_io_schedule_bits_c_bits_tag),
    .io_schedule_bits_c_bits_set(abc_mshrs_1_io_schedule_bits_c_bits_set),
    .io_schedule_bits_c_bits_way(abc_mshrs_1_io_schedule_bits_c_bits_way),
    .io_schedule_bits_c_bits_dirty(abc_mshrs_1_io_schedule_bits_c_bits_dirty),
    .io_schedule_bits_d_valid(abc_mshrs_1_io_schedule_bits_d_valid),
    .io_schedule_bits_d_bits_prio_0(abc_mshrs_1_io_schedule_bits_d_bits_prio_0),
    .io_schedule_bits_d_bits_prio_1(abc_mshrs_1_io_schedule_bits_d_bits_prio_1),
    .io_schedule_bits_d_bits_prio_2(abc_mshrs_1_io_schedule_bits_d_bits_prio_2),
    .io_schedule_bits_d_bits_control(abc_mshrs_1_io_schedule_bits_d_bits_control),
    .io_schedule_bits_d_bits_opcode(abc_mshrs_1_io_schedule_bits_d_bits_opcode),
    .io_schedule_bits_d_bits_param(abc_mshrs_1_io_schedule_bits_d_bits_param),
    .io_schedule_bits_d_bits_size(abc_mshrs_1_io_schedule_bits_d_bits_size),
    .io_schedule_bits_d_bits_source(abc_mshrs_1_io_schedule_bits_d_bits_source),
    .io_schedule_bits_d_bits_tag(abc_mshrs_1_io_schedule_bits_d_bits_tag),
    .io_schedule_bits_d_bits_offset(abc_mshrs_1_io_schedule_bits_d_bits_offset),
    .io_schedule_bits_d_bits_put(abc_mshrs_1_io_schedule_bits_d_bits_put),
    .io_schedule_bits_d_bits_set(abc_mshrs_1_io_schedule_bits_d_bits_set),
    .io_schedule_bits_d_bits_way(abc_mshrs_1_io_schedule_bits_d_bits_way),
    .io_schedule_bits_d_bits_bad(abc_mshrs_1_io_schedule_bits_d_bits_bad),
    .io_schedule_bits_e_valid(abc_mshrs_1_io_schedule_bits_e_valid),
    .io_schedule_bits_e_bits_sink(abc_mshrs_1_io_schedule_bits_e_bits_sink),
    .io_schedule_bits_x_valid(abc_mshrs_1_io_schedule_bits_x_valid),
    .io_schedule_bits_dir_valid(abc_mshrs_1_io_schedule_bits_dir_valid),
    .io_schedule_bits_dir_bits_set(abc_mshrs_1_io_schedule_bits_dir_bits_set),
    .io_schedule_bits_dir_bits_way(abc_mshrs_1_io_schedule_bits_dir_bits_way),
    .io_schedule_bits_dir_bits_data_dirty(abc_mshrs_1_io_schedule_bits_dir_bits_data_dirty),
    .io_schedule_bits_dir_bits_data_state(abc_mshrs_1_io_schedule_bits_dir_bits_data_state),
    .io_schedule_bits_dir_bits_data_clients(abc_mshrs_1_io_schedule_bits_dir_bits_data_clients),
    .io_schedule_bits_dir_bits_data_tag(abc_mshrs_1_io_schedule_bits_dir_bits_data_tag),
    .io_schedule_bits_reload(abc_mshrs_1_io_schedule_bits_reload),
    .io_sinkc_valid(abc_mshrs_1_io_sinkc_valid),
    .io_sinkc_bits_last(abc_mshrs_1_io_sinkc_bits_last),
    .io_sinkc_bits_tag(abc_mshrs_1_io_sinkc_bits_tag),
    .io_sinkc_bits_source(abc_mshrs_1_io_sinkc_bits_source),
    .io_sinkc_bits_param(abc_mshrs_1_io_sinkc_bits_param),
    .io_sinkc_bits_data(abc_mshrs_1_io_sinkc_bits_data),
    .io_sinkd_valid(abc_mshrs_1_io_sinkd_valid),
    .io_sinkd_bits_last(abc_mshrs_1_io_sinkd_bits_last),
    .io_sinkd_bits_opcode(abc_mshrs_1_io_sinkd_bits_opcode),
    .io_sinkd_bits_param(abc_mshrs_1_io_sinkd_bits_param),
    .io_sinkd_bits_sink(abc_mshrs_1_io_sinkd_bits_sink),
    .io_sinkd_bits_denied(abc_mshrs_1_io_sinkd_bits_denied),
    .io_sinke_valid(abc_mshrs_1_io_sinke_valid),
    .io_nestedwb_set(abc_mshrs_1_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshrs_1_io_nestedwb_tag),
    .io_nestedwb_b_toN(abc_mshrs_1_io_nestedwb_b_toN),
    .io_nestedwb_b_toB(abc_mshrs_1_io_nestedwb_b_toB),
    .io_nestedwb_b_clr_dirty(abc_mshrs_1_io_nestedwb_b_clr_dirty),
    .io_nestedwb_c_set_dirty(abc_mshrs_1_io_nestedwb_c_set_dirty)
  );
  MSHR abc_mshrs_2 ( // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100105.4]
    .clock(abc_mshrs_2_clock),
    .reset(abc_mshrs_2_reset),
    .io_allocate_valid(abc_mshrs_2_io_allocate_valid),
    .io_allocate_bits_prio_0(abc_mshrs_2_io_allocate_bits_prio_0),
    .io_allocate_bits_prio_1(abc_mshrs_2_io_allocate_bits_prio_1),
    .io_allocate_bits_prio_2(abc_mshrs_2_io_allocate_bits_prio_2),
    .io_allocate_bits_control(abc_mshrs_2_io_allocate_bits_control),
    .io_allocate_bits_opcode(abc_mshrs_2_io_allocate_bits_opcode),
    .io_allocate_bits_param(abc_mshrs_2_io_allocate_bits_param),
    .io_allocate_bits_size(abc_mshrs_2_io_allocate_bits_size),
    .io_allocate_bits_source(abc_mshrs_2_io_allocate_bits_source),
    .io_allocate_bits_tag(abc_mshrs_2_io_allocate_bits_tag),
    .io_allocate_bits_offset(abc_mshrs_2_io_allocate_bits_offset),
    .io_allocate_bits_put(abc_mshrs_2_io_allocate_bits_put),
    .io_allocate_bits_set(abc_mshrs_2_io_allocate_bits_set),
    .io_allocate_bits_repeat(abc_mshrs_2_io_allocate_bits_repeat),
    .io_directory_valid(abc_mshrs_2_io_directory_valid),
    .io_directory_bits_dirty(abc_mshrs_2_io_directory_bits_dirty),
    .io_directory_bits_state(abc_mshrs_2_io_directory_bits_state),
    .io_directory_bits_clients(abc_mshrs_2_io_directory_bits_clients),
    .io_directory_bits_tag(abc_mshrs_2_io_directory_bits_tag),
    .io_directory_bits_hit(abc_mshrs_2_io_directory_bits_hit),
    .io_directory_bits_way(abc_mshrs_2_io_directory_bits_way),
    .io_status_valid(abc_mshrs_2_io_status_valid),
    .io_status_bits_set(abc_mshrs_2_io_status_bits_set),
    .io_status_bits_tag(abc_mshrs_2_io_status_bits_tag),
    .io_status_bits_way(abc_mshrs_2_io_status_bits_way),
    .io_status_bits_blockB(abc_mshrs_2_io_status_bits_blockB),
    .io_status_bits_nestB(abc_mshrs_2_io_status_bits_nestB),
    .io_status_bits_blockC(abc_mshrs_2_io_status_bits_blockC),
    .io_status_bits_nestC(abc_mshrs_2_io_status_bits_nestC),
    .io_schedule_ready(abc_mshrs_2_io_schedule_ready),
    .io_schedule_valid(abc_mshrs_2_io_schedule_valid),
    .io_schedule_bits_a_valid(abc_mshrs_2_io_schedule_bits_a_valid),
    .io_schedule_bits_a_bits_tag(abc_mshrs_2_io_schedule_bits_a_bits_tag),
    .io_schedule_bits_a_bits_set(abc_mshrs_2_io_schedule_bits_a_bits_set),
    .io_schedule_bits_a_bits_param(abc_mshrs_2_io_schedule_bits_a_bits_param),
    .io_schedule_bits_a_bits_block(abc_mshrs_2_io_schedule_bits_a_bits_block),
    .io_schedule_bits_b_valid(abc_mshrs_2_io_schedule_bits_b_valid),
    .io_schedule_bits_b_bits_param(abc_mshrs_2_io_schedule_bits_b_bits_param),
    .io_schedule_bits_b_bits_tag(abc_mshrs_2_io_schedule_bits_b_bits_tag),
    .io_schedule_bits_b_bits_set(abc_mshrs_2_io_schedule_bits_b_bits_set),
    .io_schedule_bits_b_bits_clients(abc_mshrs_2_io_schedule_bits_b_bits_clients),
    .io_schedule_bits_c_valid(abc_mshrs_2_io_schedule_bits_c_valid),
    .io_schedule_bits_c_bits_opcode(abc_mshrs_2_io_schedule_bits_c_bits_opcode),
    .io_schedule_bits_c_bits_param(abc_mshrs_2_io_schedule_bits_c_bits_param),
    .io_schedule_bits_c_bits_tag(abc_mshrs_2_io_schedule_bits_c_bits_tag),
    .io_schedule_bits_c_bits_set(abc_mshrs_2_io_schedule_bits_c_bits_set),
    .io_schedule_bits_c_bits_way(abc_mshrs_2_io_schedule_bits_c_bits_way),
    .io_schedule_bits_c_bits_dirty(abc_mshrs_2_io_schedule_bits_c_bits_dirty),
    .io_schedule_bits_d_valid(abc_mshrs_2_io_schedule_bits_d_valid),
    .io_schedule_bits_d_bits_prio_0(abc_mshrs_2_io_schedule_bits_d_bits_prio_0),
    .io_schedule_bits_d_bits_prio_1(abc_mshrs_2_io_schedule_bits_d_bits_prio_1),
    .io_schedule_bits_d_bits_prio_2(abc_mshrs_2_io_schedule_bits_d_bits_prio_2),
    .io_schedule_bits_d_bits_control(abc_mshrs_2_io_schedule_bits_d_bits_control),
    .io_schedule_bits_d_bits_opcode(abc_mshrs_2_io_schedule_bits_d_bits_opcode),
    .io_schedule_bits_d_bits_param(abc_mshrs_2_io_schedule_bits_d_bits_param),
    .io_schedule_bits_d_bits_size(abc_mshrs_2_io_schedule_bits_d_bits_size),
    .io_schedule_bits_d_bits_source(abc_mshrs_2_io_schedule_bits_d_bits_source),
    .io_schedule_bits_d_bits_tag(abc_mshrs_2_io_schedule_bits_d_bits_tag),
    .io_schedule_bits_d_bits_offset(abc_mshrs_2_io_schedule_bits_d_bits_offset),
    .io_schedule_bits_d_bits_put(abc_mshrs_2_io_schedule_bits_d_bits_put),
    .io_schedule_bits_d_bits_set(abc_mshrs_2_io_schedule_bits_d_bits_set),
    .io_schedule_bits_d_bits_way(abc_mshrs_2_io_schedule_bits_d_bits_way),
    .io_schedule_bits_d_bits_bad(abc_mshrs_2_io_schedule_bits_d_bits_bad),
    .io_schedule_bits_e_valid(abc_mshrs_2_io_schedule_bits_e_valid),
    .io_schedule_bits_e_bits_sink(abc_mshrs_2_io_schedule_bits_e_bits_sink),
    .io_schedule_bits_x_valid(abc_mshrs_2_io_schedule_bits_x_valid),
    .io_schedule_bits_dir_valid(abc_mshrs_2_io_schedule_bits_dir_valid),
    .io_schedule_bits_dir_bits_set(abc_mshrs_2_io_schedule_bits_dir_bits_set),
    .io_schedule_bits_dir_bits_way(abc_mshrs_2_io_schedule_bits_dir_bits_way),
    .io_schedule_bits_dir_bits_data_dirty(abc_mshrs_2_io_schedule_bits_dir_bits_data_dirty),
    .io_schedule_bits_dir_bits_data_state(abc_mshrs_2_io_schedule_bits_dir_bits_data_state),
    .io_schedule_bits_dir_bits_data_clients(abc_mshrs_2_io_schedule_bits_dir_bits_data_clients),
    .io_schedule_bits_dir_bits_data_tag(abc_mshrs_2_io_schedule_bits_dir_bits_data_tag),
    .io_schedule_bits_reload(abc_mshrs_2_io_schedule_bits_reload),
    .io_sinkc_valid(abc_mshrs_2_io_sinkc_valid),
    .io_sinkc_bits_last(abc_mshrs_2_io_sinkc_bits_last),
    .io_sinkc_bits_tag(abc_mshrs_2_io_sinkc_bits_tag),
    .io_sinkc_bits_source(abc_mshrs_2_io_sinkc_bits_source),
    .io_sinkc_bits_param(abc_mshrs_2_io_sinkc_bits_param),
    .io_sinkc_bits_data(abc_mshrs_2_io_sinkc_bits_data),
    .io_sinkd_valid(abc_mshrs_2_io_sinkd_valid),
    .io_sinkd_bits_last(abc_mshrs_2_io_sinkd_bits_last),
    .io_sinkd_bits_opcode(abc_mshrs_2_io_sinkd_bits_opcode),
    .io_sinkd_bits_param(abc_mshrs_2_io_sinkd_bits_param),
    .io_sinkd_bits_sink(abc_mshrs_2_io_sinkd_bits_sink),
    .io_sinkd_bits_denied(abc_mshrs_2_io_sinkd_bits_denied),
    .io_sinke_valid(abc_mshrs_2_io_sinke_valid),
    .io_nestedwb_set(abc_mshrs_2_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshrs_2_io_nestedwb_tag),
    .io_nestedwb_b_toN(abc_mshrs_2_io_nestedwb_b_toN),
    .io_nestedwb_b_toB(abc_mshrs_2_io_nestedwb_b_toB),
    .io_nestedwb_b_clr_dirty(abc_mshrs_2_io_nestedwb_b_clr_dirty),
    .io_nestedwb_c_set_dirty(abc_mshrs_2_io_nestedwb_c_set_dirty)
  );
  MSHR abc_mshrs_3 ( // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100109.4]
    .clock(abc_mshrs_3_clock),
    .reset(abc_mshrs_3_reset),
    .io_allocate_valid(abc_mshrs_3_io_allocate_valid),
    .io_allocate_bits_prio_0(abc_mshrs_3_io_allocate_bits_prio_0),
    .io_allocate_bits_prio_1(abc_mshrs_3_io_allocate_bits_prio_1),
    .io_allocate_bits_prio_2(abc_mshrs_3_io_allocate_bits_prio_2),
    .io_allocate_bits_control(abc_mshrs_3_io_allocate_bits_control),
    .io_allocate_bits_opcode(abc_mshrs_3_io_allocate_bits_opcode),
    .io_allocate_bits_param(abc_mshrs_3_io_allocate_bits_param),
    .io_allocate_bits_size(abc_mshrs_3_io_allocate_bits_size),
    .io_allocate_bits_source(abc_mshrs_3_io_allocate_bits_source),
    .io_allocate_bits_tag(abc_mshrs_3_io_allocate_bits_tag),
    .io_allocate_bits_offset(abc_mshrs_3_io_allocate_bits_offset),
    .io_allocate_bits_put(abc_mshrs_3_io_allocate_bits_put),
    .io_allocate_bits_set(abc_mshrs_3_io_allocate_bits_set),
    .io_allocate_bits_repeat(abc_mshrs_3_io_allocate_bits_repeat),
    .io_directory_valid(abc_mshrs_3_io_directory_valid),
    .io_directory_bits_dirty(abc_mshrs_3_io_directory_bits_dirty),
    .io_directory_bits_state(abc_mshrs_3_io_directory_bits_state),
    .io_directory_bits_clients(abc_mshrs_3_io_directory_bits_clients),
    .io_directory_bits_tag(abc_mshrs_3_io_directory_bits_tag),
    .io_directory_bits_hit(abc_mshrs_3_io_directory_bits_hit),
    .io_directory_bits_way(abc_mshrs_3_io_directory_bits_way),
    .io_status_valid(abc_mshrs_3_io_status_valid),
    .io_status_bits_set(abc_mshrs_3_io_status_bits_set),
    .io_status_bits_tag(abc_mshrs_3_io_status_bits_tag),
    .io_status_bits_way(abc_mshrs_3_io_status_bits_way),
    .io_status_bits_blockB(abc_mshrs_3_io_status_bits_blockB),
    .io_status_bits_nestB(abc_mshrs_3_io_status_bits_nestB),
    .io_status_bits_blockC(abc_mshrs_3_io_status_bits_blockC),
    .io_status_bits_nestC(abc_mshrs_3_io_status_bits_nestC),
    .io_schedule_ready(abc_mshrs_3_io_schedule_ready),
    .io_schedule_valid(abc_mshrs_3_io_schedule_valid),
    .io_schedule_bits_a_valid(abc_mshrs_3_io_schedule_bits_a_valid),
    .io_schedule_bits_a_bits_tag(abc_mshrs_3_io_schedule_bits_a_bits_tag),
    .io_schedule_bits_a_bits_set(abc_mshrs_3_io_schedule_bits_a_bits_set),
    .io_schedule_bits_a_bits_param(abc_mshrs_3_io_schedule_bits_a_bits_param),
    .io_schedule_bits_a_bits_block(abc_mshrs_3_io_schedule_bits_a_bits_block),
    .io_schedule_bits_b_valid(abc_mshrs_3_io_schedule_bits_b_valid),
    .io_schedule_bits_b_bits_param(abc_mshrs_3_io_schedule_bits_b_bits_param),
    .io_schedule_bits_b_bits_tag(abc_mshrs_3_io_schedule_bits_b_bits_tag),
    .io_schedule_bits_b_bits_set(abc_mshrs_3_io_schedule_bits_b_bits_set),
    .io_schedule_bits_b_bits_clients(abc_mshrs_3_io_schedule_bits_b_bits_clients),
    .io_schedule_bits_c_valid(abc_mshrs_3_io_schedule_bits_c_valid),
    .io_schedule_bits_c_bits_opcode(abc_mshrs_3_io_schedule_bits_c_bits_opcode),
    .io_schedule_bits_c_bits_param(abc_mshrs_3_io_schedule_bits_c_bits_param),
    .io_schedule_bits_c_bits_tag(abc_mshrs_3_io_schedule_bits_c_bits_tag),
    .io_schedule_bits_c_bits_set(abc_mshrs_3_io_schedule_bits_c_bits_set),
    .io_schedule_bits_c_bits_way(abc_mshrs_3_io_schedule_bits_c_bits_way),
    .io_schedule_bits_c_bits_dirty(abc_mshrs_3_io_schedule_bits_c_bits_dirty),
    .io_schedule_bits_d_valid(abc_mshrs_3_io_schedule_bits_d_valid),
    .io_schedule_bits_d_bits_prio_0(abc_mshrs_3_io_schedule_bits_d_bits_prio_0),
    .io_schedule_bits_d_bits_prio_1(abc_mshrs_3_io_schedule_bits_d_bits_prio_1),
    .io_schedule_bits_d_bits_prio_2(abc_mshrs_3_io_schedule_bits_d_bits_prio_2),
    .io_schedule_bits_d_bits_control(abc_mshrs_3_io_schedule_bits_d_bits_control),
    .io_schedule_bits_d_bits_opcode(abc_mshrs_3_io_schedule_bits_d_bits_opcode),
    .io_schedule_bits_d_bits_param(abc_mshrs_3_io_schedule_bits_d_bits_param),
    .io_schedule_bits_d_bits_size(abc_mshrs_3_io_schedule_bits_d_bits_size),
    .io_schedule_bits_d_bits_source(abc_mshrs_3_io_schedule_bits_d_bits_source),
    .io_schedule_bits_d_bits_tag(abc_mshrs_3_io_schedule_bits_d_bits_tag),
    .io_schedule_bits_d_bits_offset(abc_mshrs_3_io_schedule_bits_d_bits_offset),
    .io_schedule_bits_d_bits_put(abc_mshrs_3_io_schedule_bits_d_bits_put),
    .io_schedule_bits_d_bits_set(abc_mshrs_3_io_schedule_bits_d_bits_set),
    .io_schedule_bits_d_bits_way(abc_mshrs_3_io_schedule_bits_d_bits_way),
    .io_schedule_bits_d_bits_bad(abc_mshrs_3_io_schedule_bits_d_bits_bad),
    .io_schedule_bits_e_valid(abc_mshrs_3_io_schedule_bits_e_valid),
    .io_schedule_bits_e_bits_sink(abc_mshrs_3_io_schedule_bits_e_bits_sink),
    .io_schedule_bits_x_valid(abc_mshrs_3_io_schedule_bits_x_valid),
    .io_schedule_bits_dir_valid(abc_mshrs_3_io_schedule_bits_dir_valid),
    .io_schedule_bits_dir_bits_set(abc_mshrs_3_io_schedule_bits_dir_bits_set),
    .io_schedule_bits_dir_bits_way(abc_mshrs_3_io_schedule_bits_dir_bits_way),
    .io_schedule_bits_dir_bits_data_dirty(abc_mshrs_3_io_schedule_bits_dir_bits_data_dirty),
    .io_schedule_bits_dir_bits_data_state(abc_mshrs_3_io_schedule_bits_dir_bits_data_state),
    .io_schedule_bits_dir_bits_data_clients(abc_mshrs_3_io_schedule_bits_dir_bits_data_clients),
    .io_schedule_bits_dir_bits_data_tag(abc_mshrs_3_io_schedule_bits_dir_bits_data_tag),
    .io_schedule_bits_reload(abc_mshrs_3_io_schedule_bits_reload),
    .io_sinkc_valid(abc_mshrs_3_io_sinkc_valid),
    .io_sinkc_bits_last(abc_mshrs_3_io_sinkc_bits_last),
    .io_sinkc_bits_tag(abc_mshrs_3_io_sinkc_bits_tag),
    .io_sinkc_bits_source(abc_mshrs_3_io_sinkc_bits_source),
    .io_sinkc_bits_param(abc_mshrs_3_io_sinkc_bits_param),
    .io_sinkc_bits_data(abc_mshrs_3_io_sinkc_bits_data),
    .io_sinkd_valid(abc_mshrs_3_io_sinkd_valid),
    .io_sinkd_bits_last(abc_mshrs_3_io_sinkd_bits_last),
    .io_sinkd_bits_opcode(abc_mshrs_3_io_sinkd_bits_opcode),
    .io_sinkd_bits_param(abc_mshrs_3_io_sinkd_bits_param),
    .io_sinkd_bits_sink(abc_mshrs_3_io_sinkd_bits_sink),
    .io_sinkd_bits_denied(abc_mshrs_3_io_sinkd_bits_denied),
    .io_sinke_valid(abc_mshrs_3_io_sinke_valid),
    .io_nestedwb_set(abc_mshrs_3_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshrs_3_io_nestedwb_tag),
    .io_nestedwb_b_toN(abc_mshrs_3_io_nestedwb_b_toN),
    .io_nestedwb_b_toB(abc_mshrs_3_io_nestedwb_b_toB),
    .io_nestedwb_b_clr_dirty(abc_mshrs_3_io_nestedwb_b_clr_dirty),
    .io_nestedwb_c_set_dirty(abc_mshrs_3_io_nestedwb_c_set_dirty)
  );
  MSHR abc_mshrs_4 ( // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100113.4]
    .clock(abc_mshrs_4_clock),
    .reset(abc_mshrs_4_reset),
    .io_allocate_valid(abc_mshrs_4_io_allocate_valid),
    .io_allocate_bits_prio_0(abc_mshrs_4_io_allocate_bits_prio_0),
    .io_allocate_bits_prio_1(abc_mshrs_4_io_allocate_bits_prio_1),
    .io_allocate_bits_prio_2(abc_mshrs_4_io_allocate_bits_prio_2),
    .io_allocate_bits_control(abc_mshrs_4_io_allocate_bits_control),
    .io_allocate_bits_opcode(abc_mshrs_4_io_allocate_bits_opcode),
    .io_allocate_bits_param(abc_mshrs_4_io_allocate_bits_param),
    .io_allocate_bits_size(abc_mshrs_4_io_allocate_bits_size),
    .io_allocate_bits_source(abc_mshrs_4_io_allocate_bits_source),
    .io_allocate_bits_tag(abc_mshrs_4_io_allocate_bits_tag),
    .io_allocate_bits_offset(abc_mshrs_4_io_allocate_bits_offset),
    .io_allocate_bits_put(abc_mshrs_4_io_allocate_bits_put),
    .io_allocate_bits_set(abc_mshrs_4_io_allocate_bits_set),
    .io_allocate_bits_repeat(abc_mshrs_4_io_allocate_bits_repeat),
    .io_directory_valid(abc_mshrs_4_io_directory_valid),
    .io_directory_bits_dirty(abc_mshrs_4_io_directory_bits_dirty),
    .io_directory_bits_state(abc_mshrs_4_io_directory_bits_state),
    .io_directory_bits_clients(abc_mshrs_4_io_directory_bits_clients),
    .io_directory_bits_tag(abc_mshrs_4_io_directory_bits_tag),
    .io_directory_bits_hit(abc_mshrs_4_io_directory_bits_hit),
    .io_directory_bits_way(abc_mshrs_4_io_directory_bits_way),
    .io_status_valid(abc_mshrs_4_io_status_valid),
    .io_status_bits_set(abc_mshrs_4_io_status_bits_set),
    .io_status_bits_tag(abc_mshrs_4_io_status_bits_tag),
    .io_status_bits_way(abc_mshrs_4_io_status_bits_way),
    .io_status_bits_blockB(abc_mshrs_4_io_status_bits_blockB),
    .io_status_bits_nestB(abc_mshrs_4_io_status_bits_nestB),
    .io_status_bits_blockC(abc_mshrs_4_io_status_bits_blockC),
    .io_status_bits_nestC(abc_mshrs_4_io_status_bits_nestC),
    .io_schedule_ready(abc_mshrs_4_io_schedule_ready),
    .io_schedule_valid(abc_mshrs_4_io_schedule_valid),
    .io_schedule_bits_a_valid(abc_mshrs_4_io_schedule_bits_a_valid),
    .io_schedule_bits_a_bits_tag(abc_mshrs_4_io_schedule_bits_a_bits_tag),
    .io_schedule_bits_a_bits_set(abc_mshrs_4_io_schedule_bits_a_bits_set),
    .io_schedule_bits_a_bits_param(abc_mshrs_4_io_schedule_bits_a_bits_param),
    .io_schedule_bits_a_bits_block(abc_mshrs_4_io_schedule_bits_a_bits_block),
    .io_schedule_bits_b_valid(abc_mshrs_4_io_schedule_bits_b_valid),
    .io_schedule_bits_b_bits_param(abc_mshrs_4_io_schedule_bits_b_bits_param),
    .io_schedule_bits_b_bits_tag(abc_mshrs_4_io_schedule_bits_b_bits_tag),
    .io_schedule_bits_b_bits_set(abc_mshrs_4_io_schedule_bits_b_bits_set),
    .io_schedule_bits_b_bits_clients(abc_mshrs_4_io_schedule_bits_b_bits_clients),
    .io_schedule_bits_c_valid(abc_mshrs_4_io_schedule_bits_c_valid),
    .io_schedule_bits_c_bits_opcode(abc_mshrs_4_io_schedule_bits_c_bits_opcode),
    .io_schedule_bits_c_bits_param(abc_mshrs_4_io_schedule_bits_c_bits_param),
    .io_schedule_bits_c_bits_tag(abc_mshrs_4_io_schedule_bits_c_bits_tag),
    .io_schedule_bits_c_bits_set(abc_mshrs_4_io_schedule_bits_c_bits_set),
    .io_schedule_bits_c_bits_way(abc_mshrs_4_io_schedule_bits_c_bits_way),
    .io_schedule_bits_c_bits_dirty(abc_mshrs_4_io_schedule_bits_c_bits_dirty),
    .io_schedule_bits_d_valid(abc_mshrs_4_io_schedule_bits_d_valid),
    .io_schedule_bits_d_bits_prio_0(abc_mshrs_4_io_schedule_bits_d_bits_prio_0),
    .io_schedule_bits_d_bits_prio_1(abc_mshrs_4_io_schedule_bits_d_bits_prio_1),
    .io_schedule_bits_d_bits_prio_2(abc_mshrs_4_io_schedule_bits_d_bits_prio_2),
    .io_schedule_bits_d_bits_control(abc_mshrs_4_io_schedule_bits_d_bits_control),
    .io_schedule_bits_d_bits_opcode(abc_mshrs_4_io_schedule_bits_d_bits_opcode),
    .io_schedule_bits_d_bits_param(abc_mshrs_4_io_schedule_bits_d_bits_param),
    .io_schedule_bits_d_bits_size(abc_mshrs_4_io_schedule_bits_d_bits_size),
    .io_schedule_bits_d_bits_source(abc_mshrs_4_io_schedule_bits_d_bits_source),
    .io_schedule_bits_d_bits_tag(abc_mshrs_4_io_schedule_bits_d_bits_tag),
    .io_schedule_bits_d_bits_offset(abc_mshrs_4_io_schedule_bits_d_bits_offset),
    .io_schedule_bits_d_bits_put(abc_mshrs_4_io_schedule_bits_d_bits_put),
    .io_schedule_bits_d_bits_set(abc_mshrs_4_io_schedule_bits_d_bits_set),
    .io_schedule_bits_d_bits_way(abc_mshrs_4_io_schedule_bits_d_bits_way),
    .io_schedule_bits_d_bits_bad(abc_mshrs_4_io_schedule_bits_d_bits_bad),
    .io_schedule_bits_e_valid(abc_mshrs_4_io_schedule_bits_e_valid),
    .io_schedule_bits_e_bits_sink(abc_mshrs_4_io_schedule_bits_e_bits_sink),
    .io_schedule_bits_x_valid(abc_mshrs_4_io_schedule_bits_x_valid),
    .io_schedule_bits_dir_valid(abc_mshrs_4_io_schedule_bits_dir_valid),
    .io_schedule_bits_dir_bits_set(abc_mshrs_4_io_schedule_bits_dir_bits_set),
    .io_schedule_bits_dir_bits_way(abc_mshrs_4_io_schedule_bits_dir_bits_way),
    .io_schedule_bits_dir_bits_data_dirty(abc_mshrs_4_io_schedule_bits_dir_bits_data_dirty),
    .io_schedule_bits_dir_bits_data_state(abc_mshrs_4_io_schedule_bits_dir_bits_data_state),
    .io_schedule_bits_dir_bits_data_clients(abc_mshrs_4_io_schedule_bits_dir_bits_data_clients),
    .io_schedule_bits_dir_bits_data_tag(abc_mshrs_4_io_schedule_bits_dir_bits_data_tag),
    .io_schedule_bits_reload(abc_mshrs_4_io_schedule_bits_reload),
    .io_sinkc_valid(abc_mshrs_4_io_sinkc_valid),
    .io_sinkc_bits_last(abc_mshrs_4_io_sinkc_bits_last),
    .io_sinkc_bits_tag(abc_mshrs_4_io_sinkc_bits_tag),
    .io_sinkc_bits_source(abc_mshrs_4_io_sinkc_bits_source),
    .io_sinkc_bits_param(abc_mshrs_4_io_sinkc_bits_param),
    .io_sinkc_bits_data(abc_mshrs_4_io_sinkc_bits_data),
    .io_sinkd_valid(abc_mshrs_4_io_sinkd_valid),
    .io_sinkd_bits_last(abc_mshrs_4_io_sinkd_bits_last),
    .io_sinkd_bits_opcode(abc_mshrs_4_io_sinkd_bits_opcode),
    .io_sinkd_bits_param(abc_mshrs_4_io_sinkd_bits_param),
    .io_sinkd_bits_sink(abc_mshrs_4_io_sinkd_bits_sink),
    .io_sinkd_bits_denied(abc_mshrs_4_io_sinkd_bits_denied),
    .io_sinke_valid(abc_mshrs_4_io_sinke_valid),
    .io_nestedwb_set(abc_mshrs_4_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshrs_4_io_nestedwb_tag),
    .io_nestedwb_b_toN(abc_mshrs_4_io_nestedwb_b_toN),
    .io_nestedwb_b_toB(abc_mshrs_4_io_nestedwb_b_toB),
    .io_nestedwb_b_clr_dirty(abc_mshrs_4_io_nestedwb_b_clr_dirty),
    .io_nestedwb_c_set_dirty(abc_mshrs_4_io_nestedwb_c_set_dirty)
  );
  MSHR bc_mshr ( // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100117.4]
    .clock(bc_mshr_clock),
    .reset(bc_mshr_reset),
    .io_allocate_valid(bc_mshr_io_allocate_valid),
    .io_allocate_bits_prio_0(bc_mshr_io_allocate_bits_prio_0),
    .io_allocate_bits_prio_1(bc_mshr_io_allocate_bits_prio_1),
    .io_allocate_bits_prio_2(bc_mshr_io_allocate_bits_prio_2),
    .io_allocate_bits_control(bc_mshr_io_allocate_bits_control),
    .io_allocate_bits_opcode(bc_mshr_io_allocate_bits_opcode),
    .io_allocate_bits_param(bc_mshr_io_allocate_bits_param),
    .io_allocate_bits_size(bc_mshr_io_allocate_bits_size),
    .io_allocate_bits_source(bc_mshr_io_allocate_bits_source),
    .io_allocate_bits_tag(bc_mshr_io_allocate_bits_tag),
    .io_allocate_bits_offset(bc_mshr_io_allocate_bits_offset),
    .io_allocate_bits_put(bc_mshr_io_allocate_bits_put),
    .io_allocate_bits_set(bc_mshr_io_allocate_bits_set),
    .io_allocate_bits_repeat(bc_mshr_io_allocate_bits_repeat),
    .io_directory_valid(bc_mshr_io_directory_valid),
    .io_directory_bits_dirty(bc_mshr_io_directory_bits_dirty),
    .io_directory_bits_state(bc_mshr_io_directory_bits_state),
    .io_directory_bits_clients(bc_mshr_io_directory_bits_clients),
    .io_directory_bits_tag(bc_mshr_io_directory_bits_tag),
    .io_directory_bits_hit(bc_mshr_io_directory_bits_hit),
    .io_directory_bits_way(bc_mshr_io_directory_bits_way),
    .io_status_valid(bc_mshr_io_status_valid),
    .io_status_bits_set(bc_mshr_io_status_bits_set),
    .io_status_bits_tag(bc_mshr_io_status_bits_tag),
    .io_status_bits_way(bc_mshr_io_status_bits_way),
    .io_status_bits_blockB(bc_mshr_io_status_bits_blockB),
    .io_status_bits_nestB(bc_mshr_io_status_bits_nestB),
    .io_status_bits_blockC(bc_mshr_io_status_bits_blockC),
    .io_status_bits_nestC(bc_mshr_io_status_bits_nestC),
    .io_schedule_ready(bc_mshr_io_schedule_ready),
    .io_schedule_valid(bc_mshr_io_schedule_valid),
    .io_schedule_bits_a_valid(bc_mshr_io_schedule_bits_a_valid),
    .io_schedule_bits_a_bits_tag(bc_mshr_io_schedule_bits_a_bits_tag),
    .io_schedule_bits_a_bits_set(bc_mshr_io_schedule_bits_a_bits_set),
    .io_schedule_bits_a_bits_param(bc_mshr_io_schedule_bits_a_bits_param),
    .io_schedule_bits_a_bits_block(bc_mshr_io_schedule_bits_a_bits_block),
    .io_schedule_bits_b_valid(bc_mshr_io_schedule_bits_b_valid),
    .io_schedule_bits_b_bits_param(bc_mshr_io_schedule_bits_b_bits_param),
    .io_schedule_bits_b_bits_tag(bc_mshr_io_schedule_bits_b_bits_tag),
    .io_schedule_bits_b_bits_set(bc_mshr_io_schedule_bits_b_bits_set),
    .io_schedule_bits_b_bits_clients(bc_mshr_io_schedule_bits_b_bits_clients),
    .io_schedule_bits_c_valid(bc_mshr_io_schedule_bits_c_valid),
    .io_schedule_bits_c_bits_opcode(bc_mshr_io_schedule_bits_c_bits_opcode),
    .io_schedule_bits_c_bits_param(bc_mshr_io_schedule_bits_c_bits_param),
    .io_schedule_bits_c_bits_tag(bc_mshr_io_schedule_bits_c_bits_tag),
    .io_schedule_bits_c_bits_set(bc_mshr_io_schedule_bits_c_bits_set),
    .io_schedule_bits_c_bits_way(bc_mshr_io_schedule_bits_c_bits_way),
    .io_schedule_bits_c_bits_dirty(bc_mshr_io_schedule_bits_c_bits_dirty),
    .io_schedule_bits_d_valid(bc_mshr_io_schedule_bits_d_valid),
    .io_schedule_bits_d_bits_prio_0(bc_mshr_io_schedule_bits_d_bits_prio_0),
    .io_schedule_bits_d_bits_prio_1(bc_mshr_io_schedule_bits_d_bits_prio_1),
    .io_schedule_bits_d_bits_prio_2(bc_mshr_io_schedule_bits_d_bits_prio_2),
    .io_schedule_bits_d_bits_control(bc_mshr_io_schedule_bits_d_bits_control),
    .io_schedule_bits_d_bits_opcode(bc_mshr_io_schedule_bits_d_bits_opcode),
    .io_schedule_bits_d_bits_param(bc_mshr_io_schedule_bits_d_bits_param),
    .io_schedule_bits_d_bits_size(bc_mshr_io_schedule_bits_d_bits_size),
    .io_schedule_bits_d_bits_source(bc_mshr_io_schedule_bits_d_bits_source),
    .io_schedule_bits_d_bits_tag(bc_mshr_io_schedule_bits_d_bits_tag),
    .io_schedule_bits_d_bits_offset(bc_mshr_io_schedule_bits_d_bits_offset),
    .io_schedule_bits_d_bits_put(bc_mshr_io_schedule_bits_d_bits_put),
    .io_schedule_bits_d_bits_set(bc_mshr_io_schedule_bits_d_bits_set),
    .io_schedule_bits_d_bits_way(bc_mshr_io_schedule_bits_d_bits_way),
    .io_schedule_bits_d_bits_bad(bc_mshr_io_schedule_bits_d_bits_bad),
    .io_schedule_bits_e_valid(bc_mshr_io_schedule_bits_e_valid),
    .io_schedule_bits_e_bits_sink(bc_mshr_io_schedule_bits_e_bits_sink),
    .io_schedule_bits_x_valid(bc_mshr_io_schedule_bits_x_valid),
    .io_schedule_bits_dir_valid(bc_mshr_io_schedule_bits_dir_valid),
    .io_schedule_bits_dir_bits_set(bc_mshr_io_schedule_bits_dir_bits_set),
    .io_schedule_bits_dir_bits_way(bc_mshr_io_schedule_bits_dir_bits_way),
    .io_schedule_bits_dir_bits_data_dirty(bc_mshr_io_schedule_bits_dir_bits_data_dirty),
    .io_schedule_bits_dir_bits_data_state(bc_mshr_io_schedule_bits_dir_bits_data_state),
    .io_schedule_bits_dir_bits_data_clients(bc_mshr_io_schedule_bits_dir_bits_data_clients),
    .io_schedule_bits_dir_bits_data_tag(bc_mshr_io_schedule_bits_dir_bits_data_tag),
    .io_schedule_bits_reload(bc_mshr_io_schedule_bits_reload),
    .io_sinkc_valid(bc_mshr_io_sinkc_valid),
    .io_sinkc_bits_last(bc_mshr_io_sinkc_bits_last),
    .io_sinkc_bits_tag(bc_mshr_io_sinkc_bits_tag),
    .io_sinkc_bits_source(bc_mshr_io_sinkc_bits_source),
    .io_sinkc_bits_param(bc_mshr_io_sinkc_bits_param),
    .io_sinkc_bits_data(bc_mshr_io_sinkc_bits_data),
    .io_sinkd_valid(bc_mshr_io_sinkd_valid),
    .io_sinkd_bits_last(bc_mshr_io_sinkd_bits_last),
    .io_sinkd_bits_opcode(bc_mshr_io_sinkd_bits_opcode),
    .io_sinkd_bits_param(bc_mshr_io_sinkd_bits_param),
    .io_sinkd_bits_sink(bc_mshr_io_sinkd_bits_sink),
    .io_sinkd_bits_denied(bc_mshr_io_sinkd_bits_denied),
    .io_sinke_valid(bc_mshr_io_sinke_valid),
    .io_nestedwb_set(bc_mshr_io_nestedwb_set),
    .io_nestedwb_tag(bc_mshr_io_nestedwb_tag),
    .io_nestedwb_b_toN(bc_mshr_io_nestedwb_b_toN),
    .io_nestedwb_b_toB(bc_mshr_io_nestedwb_b_toB),
    .io_nestedwb_b_clr_dirty(bc_mshr_io_nestedwb_b_clr_dirty),
    .io_nestedwb_c_set_dirty(bc_mshr_io_nestedwb_c_set_dirty)
  );
  MSHR c_mshr ( // @[Scheduler.scala 69:46:chipyard.TestHarness.RocketConfig.fir@100121.4]
    .clock(c_mshr_clock),
    .reset(c_mshr_reset),
    .io_allocate_valid(c_mshr_io_allocate_valid),
    .io_allocate_bits_prio_0(c_mshr_io_allocate_bits_prio_0),
    .io_allocate_bits_prio_1(c_mshr_io_allocate_bits_prio_1),
    .io_allocate_bits_prio_2(c_mshr_io_allocate_bits_prio_2),
    .io_allocate_bits_control(c_mshr_io_allocate_bits_control),
    .io_allocate_bits_opcode(c_mshr_io_allocate_bits_opcode),
    .io_allocate_bits_param(c_mshr_io_allocate_bits_param),
    .io_allocate_bits_size(c_mshr_io_allocate_bits_size),
    .io_allocate_bits_source(c_mshr_io_allocate_bits_source),
    .io_allocate_bits_tag(c_mshr_io_allocate_bits_tag),
    .io_allocate_bits_offset(c_mshr_io_allocate_bits_offset),
    .io_allocate_bits_put(c_mshr_io_allocate_bits_put),
    .io_allocate_bits_set(c_mshr_io_allocate_bits_set),
    .io_allocate_bits_repeat(c_mshr_io_allocate_bits_repeat),
    .io_directory_valid(c_mshr_io_directory_valid),
    .io_directory_bits_dirty(c_mshr_io_directory_bits_dirty),
    .io_directory_bits_state(c_mshr_io_directory_bits_state),
    .io_directory_bits_clients(c_mshr_io_directory_bits_clients),
    .io_directory_bits_tag(c_mshr_io_directory_bits_tag),
    .io_directory_bits_hit(c_mshr_io_directory_bits_hit),
    .io_directory_bits_way(c_mshr_io_directory_bits_way),
    .io_status_valid(c_mshr_io_status_valid),
    .io_status_bits_set(c_mshr_io_status_bits_set),
    .io_status_bits_tag(c_mshr_io_status_bits_tag),
    .io_status_bits_way(c_mshr_io_status_bits_way),
    .io_status_bits_blockB(c_mshr_io_status_bits_blockB),
    .io_status_bits_nestB(c_mshr_io_status_bits_nestB),
    .io_status_bits_blockC(c_mshr_io_status_bits_blockC),
    .io_status_bits_nestC(c_mshr_io_status_bits_nestC),
    .io_schedule_ready(c_mshr_io_schedule_ready),
    .io_schedule_valid(c_mshr_io_schedule_valid),
    .io_schedule_bits_a_valid(c_mshr_io_schedule_bits_a_valid),
    .io_schedule_bits_a_bits_tag(c_mshr_io_schedule_bits_a_bits_tag),
    .io_schedule_bits_a_bits_set(c_mshr_io_schedule_bits_a_bits_set),
    .io_schedule_bits_a_bits_param(c_mshr_io_schedule_bits_a_bits_param),
    .io_schedule_bits_a_bits_block(c_mshr_io_schedule_bits_a_bits_block),
    .io_schedule_bits_b_valid(c_mshr_io_schedule_bits_b_valid),
    .io_schedule_bits_b_bits_param(c_mshr_io_schedule_bits_b_bits_param),
    .io_schedule_bits_b_bits_tag(c_mshr_io_schedule_bits_b_bits_tag),
    .io_schedule_bits_b_bits_set(c_mshr_io_schedule_bits_b_bits_set),
    .io_schedule_bits_b_bits_clients(c_mshr_io_schedule_bits_b_bits_clients),
    .io_schedule_bits_c_valid(c_mshr_io_schedule_bits_c_valid),
    .io_schedule_bits_c_bits_opcode(c_mshr_io_schedule_bits_c_bits_opcode),
    .io_schedule_bits_c_bits_param(c_mshr_io_schedule_bits_c_bits_param),
    .io_schedule_bits_c_bits_tag(c_mshr_io_schedule_bits_c_bits_tag),
    .io_schedule_bits_c_bits_set(c_mshr_io_schedule_bits_c_bits_set),
    .io_schedule_bits_c_bits_way(c_mshr_io_schedule_bits_c_bits_way),
    .io_schedule_bits_c_bits_dirty(c_mshr_io_schedule_bits_c_bits_dirty),
    .io_schedule_bits_d_valid(c_mshr_io_schedule_bits_d_valid),
    .io_schedule_bits_d_bits_prio_0(c_mshr_io_schedule_bits_d_bits_prio_0),
    .io_schedule_bits_d_bits_prio_1(c_mshr_io_schedule_bits_d_bits_prio_1),
    .io_schedule_bits_d_bits_prio_2(c_mshr_io_schedule_bits_d_bits_prio_2),
    .io_schedule_bits_d_bits_control(c_mshr_io_schedule_bits_d_bits_control),
    .io_schedule_bits_d_bits_opcode(c_mshr_io_schedule_bits_d_bits_opcode),
    .io_schedule_bits_d_bits_param(c_mshr_io_schedule_bits_d_bits_param),
    .io_schedule_bits_d_bits_size(c_mshr_io_schedule_bits_d_bits_size),
    .io_schedule_bits_d_bits_source(c_mshr_io_schedule_bits_d_bits_source),
    .io_schedule_bits_d_bits_tag(c_mshr_io_schedule_bits_d_bits_tag),
    .io_schedule_bits_d_bits_offset(c_mshr_io_schedule_bits_d_bits_offset),
    .io_schedule_bits_d_bits_put(c_mshr_io_schedule_bits_d_bits_put),
    .io_schedule_bits_d_bits_set(c_mshr_io_schedule_bits_d_bits_set),
    .io_schedule_bits_d_bits_way(c_mshr_io_schedule_bits_d_bits_way),
    .io_schedule_bits_d_bits_bad(c_mshr_io_schedule_bits_d_bits_bad),
    .io_schedule_bits_e_valid(c_mshr_io_schedule_bits_e_valid),
    .io_schedule_bits_e_bits_sink(c_mshr_io_schedule_bits_e_bits_sink),
    .io_schedule_bits_x_valid(c_mshr_io_schedule_bits_x_valid),
    .io_schedule_bits_dir_valid(c_mshr_io_schedule_bits_dir_valid),
    .io_schedule_bits_dir_bits_set(c_mshr_io_schedule_bits_dir_bits_set),
    .io_schedule_bits_dir_bits_way(c_mshr_io_schedule_bits_dir_bits_way),
    .io_schedule_bits_dir_bits_data_dirty(c_mshr_io_schedule_bits_dir_bits_data_dirty),
    .io_schedule_bits_dir_bits_data_state(c_mshr_io_schedule_bits_dir_bits_data_state),
    .io_schedule_bits_dir_bits_data_clients(c_mshr_io_schedule_bits_dir_bits_data_clients),
    .io_schedule_bits_dir_bits_data_tag(c_mshr_io_schedule_bits_dir_bits_data_tag),
    .io_schedule_bits_reload(c_mshr_io_schedule_bits_reload),
    .io_sinkc_valid(c_mshr_io_sinkc_valid),
    .io_sinkc_bits_last(c_mshr_io_sinkc_bits_last),
    .io_sinkc_bits_tag(c_mshr_io_sinkc_bits_tag),
    .io_sinkc_bits_source(c_mshr_io_sinkc_bits_source),
    .io_sinkc_bits_param(c_mshr_io_sinkc_bits_param),
    .io_sinkc_bits_data(c_mshr_io_sinkc_bits_data),
    .io_sinkd_valid(c_mshr_io_sinkd_valid),
    .io_sinkd_bits_last(c_mshr_io_sinkd_bits_last),
    .io_sinkd_bits_opcode(c_mshr_io_sinkd_bits_opcode),
    .io_sinkd_bits_param(c_mshr_io_sinkd_bits_param),
    .io_sinkd_bits_sink(c_mshr_io_sinkd_bits_sink),
    .io_sinkd_bits_denied(c_mshr_io_sinkd_bits_denied),
    .io_sinke_valid(c_mshr_io_sinke_valid),
    .io_nestedwb_set(c_mshr_io_nestedwb_set),
    .io_nestedwb_tag(c_mshr_io_nestedwb_tag),
    .io_nestedwb_b_toN(c_mshr_io_nestedwb_b_toN),
    .io_nestedwb_b_toB(c_mshr_io_nestedwb_b_toB),
    .io_nestedwb_b_clr_dirty(c_mshr_io_nestedwb_b_clr_dirty),
    .io_nestedwb_c_set_dirty(c_mshr_io_nestedwb_c_set_dirty)
  );
  assign _T = sinkC_io_resp_bits_set == abc_mshrs_0_io_status_bits_set; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100127.4]
  assign _T_2 = sinkD_io_resp_bits_source == 3'h0; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100130.4]
  assign _T_4 = sinkE_io_resp_bits_sink == 3'h0; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100133.4]
  assign _T_6 = sinkC_io_resp_bits_set == abc_mshrs_1_io_status_bits_set; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100140.4]
  assign _T_8 = sinkD_io_resp_bits_source == 3'h1; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100143.4]
  assign _T_10 = sinkE_io_resp_bits_sink == 3'h1; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100146.4]
  assign _T_12 = sinkC_io_resp_bits_set == abc_mshrs_2_io_status_bits_set; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100153.4]
  assign _T_14 = sinkD_io_resp_bits_source == 3'h2; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100156.4]
  assign _T_16 = sinkE_io_resp_bits_sink == 3'h2; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100159.4]
  assign _T_18 = sinkC_io_resp_bits_set == abc_mshrs_3_io_status_bits_set; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100166.4]
  assign _T_20 = sinkD_io_resp_bits_source == 3'h3; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100169.4]
  assign _T_22 = sinkE_io_resp_bits_sink == 3'h3; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100172.4]
  assign _T_24 = sinkC_io_resp_bits_set == abc_mshrs_4_io_status_bits_set; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100179.4]
  assign _T_26 = sinkD_io_resp_bits_source == 3'h4; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100182.4]
  assign _T_28 = sinkE_io_resp_bits_sink == 3'h4; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100185.4]
  assign _T_30 = sinkC_io_resp_bits_set == bc_mshr_io_status_bits_set; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100192.4]
  assign _T_32 = sinkD_io_resp_bits_source == 3'h5; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100195.4]
  assign _T_34 = sinkE_io_resp_bits_sink == 3'h5; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100198.4]
  assign _T_36 = sinkC_io_resp_bits_set == c_mshr_io_status_bits_set; // @[Scheduler.scala 77:71:chipyard.TestHarness.RocketConfig.fir@100205.4]
  assign _T_38 = sinkD_io_resp_bits_source == 3'h6; // @[Scheduler.scala 78:74:chipyard.TestHarness.RocketConfig.fir@100208.4]
  assign _T_40 = sinkE_io_resp_bits_sink == 3'h6; // @[Scheduler.scala 79:74:chipyard.TestHarness.RocketConfig.fir@100211.4]
  assign _T_42 = abc_mshrs_0_io_status_bits_set == bc_mshr_io_status_bits_set; // @[Scheduler.scala 88:54:chipyard.TestHarness.RocketConfig.fir@100218.4]
  assign _T_43 = bc_mshr_io_status_valid & _T_42; // @[Scheduler.scala 88:30:chipyard.TestHarness.RocketConfig.fir@100219.4]
  assign _T_44 = abc_mshrs_0_io_status_bits_set == c_mshr_io_status_bits_set; // @[Scheduler.scala 89:54:chipyard.TestHarness.RocketConfig.fir@100220.4]
  assign _T_45 = c_mshr_io_status_valid & _T_44; // @[Scheduler.scala 89:30:chipyard.TestHarness.RocketConfig.fir@100221.4]
  assign mshr_stall_0 = _T_43 | _T_45; // @[Scheduler.scala 88:86:chipyard.TestHarness.RocketConfig.fir@100222.4]
  assign _T_46 = abc_mshrs_1_io_status_bits_set == bc_mshr_io_status_bits_set; // @[Scheduler.scala 88:54:chipyard.TestHarness.RocketConfig.fir@100223.4]
  assign _T_47 = bc_mshr_io_status_valid & _T_46; // @[Scheduler.scala 88:30:chipyard.TestHarness.RocketConfig.fir@100224.4]
  assign _T_48 = abc_mshrs_1_io_status_bits_set == c_mshr_io_status_bits_set; // @[Scheduler.scala 89:54:chipyard.TestHarness.RocketConfig.fir@100225.4]
  assign _T_49 = c_mshr_io_status_valid & _T_48; // @[Scheduler.scala 89:30:chipyard.TestHarness.RocketConfig.fir@100226.4]
  assign mshr_stall_1 = _T_47 | _T_49; // @[Scheduler.scala 88:86:chipyard.TestHarness.RocketConfig.fir@100227.4]
  assign _T_50 = abc_mshrs_2_io_status_bits_set == bc_mshr_io_status_bits_set; // @[Scheduler.scala 88:54:chipyard.TestHarness.RocketConfig.fir@100228.4]
  assign _T_51 = bc_mshr_io_status_valid & _T_50; // @[Scheduler.scala 88:30:chipyard.TestHarness.RocketConfig.fir@100229.4]
  assign _T_52 = abc_mshrs_2_io_status_bits_set == c_mshr_io_status_bits_set; // @[Scheduler.scala 89:54:chipyard.TestHarness.RocketConfig.fir@100230.4]
  assign _T_53 = c_mshr_io_status_valid & _T_52; // @[Scheduler.scala 89:30:chipyard.TestHarness.RocketConfig.fir@100231.4]
  assign mshr_stall_2 = _T_51 | _T_53; // @[Scheduler.scala 88:86:chipyard.TestHarness.RocketConfig.fir@100232.4]
  assign _T_54 = abc_mshrs_3_io_status_bits_set == bc_mshr_io_status_bits_set; // @[Scheduler.scala 88:54:chipyard.TestHarness.RocketConfig.fir@100233.4]
  assign _T_55 = bc_mshr_io_status_valid & _T_54; // @[Scheduler.scala 88:30:chipyard.TestHarness.RocketConfig.fir@100234.4]
  assign _T_56 = abc_mshrs_3_io_status_bits_set == c_mshr_io_status_bits_set; // @[Scheduler.scala 89:54:chipyard.TestHarness.RocketConfig.fir@100235.4]
  assign _T_57 = c_mshr_io_status_valid & _T_56; // @[Scheduler.scala 89:30:chipyard.TestHarness.RocketConfig.fir@100236.4]
  assign mshr_stall_3 = _T_55 | _T_57; // @[Scheduler.scala 88:86:chipyard.TestHarness.RocketConfig.fir@100237.4]
  assign _T_58 = abc_mshrs_4_io_status_bits_set == bc_mshr_io_status_bits_set; // @[Scheduler.scala 88:54:chipyard.TestHarness.RocketConfig.fir@100238.4]
  assign _T_59 = bc_mshr_io_status_valid & _T_58; // @[Scheduler.scala 88:30:chipyard.TestHarness.RocketConfig.fir@100239.4]
  assign _T_60 = abc_mshrs_4_io_status_bits_set == c_mshr_io_status_bits_set; // @[Scheduler.scala 89:54:chipyard.TestHarness.RocketConfig.fir@100240.4]
  assign _T_61 = c_mshr_io_status_valid & _T_60; // @[Scheduler.scala 89:30:chipyard.TestHarness.RocketConfig.fir@100241.4]
  assign mshr_stall_4 = _T_59 | _T_61; // @[Scheduler.scala 88:86:chipyard.TestHarness.RocketConfig.fir@100242.4]
  assign _T_62 = bc_mshr_io_status_bits_set == c_mshr_io_status_bits_set; // @[Scheduler.scala 92:58:chipyard.TestHarness.RocketConfig.fir@100243.4]
  assign mshr_stall_5 = c_mshr_io_status_valid & _T_62; // @[Scheduler.scala 92:28:chipyard.TestHarness.RocketConfig.fir@100244.4]
  assign _T_67 = ~mshr_stall_0; // @[Scheduler.scala 105:28:chipyard.TestHarness.RocketConfig.fir@100254.4]
  assign _T_68 = abc_mshrs_0_io_schedule_valid & _T_67; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100255.4]
  assign _T_69 = ~abc_mshrs_0_io_schedule_bits_a_valid; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100256.4]
  assign _T_70 = sourceA_io_req_ready | _T_69; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100257.4]
  assign _T_71 = _T_68 & _T_70; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100258.4]
  assign _T_72 = ~abc_mshrs_0_io_schedule_bits_b_valid; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100259.4]
  assign _T_73 = sourceB_io_req_ready | _T_72; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100260.4]
  assign _T_74 = _T_71 & _T_73; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100261.4]
  assign _T_75 = ~abc_mshrs_0_io_schedule_bits_c_valid; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100262.4]
  assign _T_76 = sourceC_io_req_ready | _T_75; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100263.4]
  assign _T_77 = _T_74 & _T_76; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100264.4]
  assign _T_78 = ~abc_mshrs_0_io_schedule_bits_d_valid; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100265.4]
  assign _T_79 = sourceD_io_req_ready | _T_78; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100266.4]
  assign _T_80 = _T_77 & _T_79; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100267.4]
  assign _T_81 = ~abc_mshrs_0_io_schedule_bits_e_valid; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100268.4]
  assign _T_82 = sourceE_io_req_ready | _T_81; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100269.4]
  assign _T_83 = _T_80 & _T_82; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100270.4]
  assign _T_84 = ~abc_mshrs_0_io_schedule_bits_x_valid; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100271.4]
  assign _T_85 = sourceX_io_req_ready | _T_84; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100272.4]
  assign _T_86 = _T_83 & _T_85; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100273.4]
  assign _T_87 = ~abc_mshrs_0_io_schedule_bits_dir_valid; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100274.4]
  assign _T_88 = directory_io_write_ready | _T_87; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100275.4]
  assign _T_89 = _T_86 & _T_88; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100276.4]
  assign _T_90 = ~mshr_stall_1; // @[Scheduler.scala 105:28:chipyard.TestHarness.RocketConfig.fir@100277.4]
  assign _T_91 = abc_mshrs_1_io_schedule_valid & _T_90; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100278.4]
  assign _T_92 = ~abc_mshrs_1_io_schedule_bits_a_valid; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100279.4]
  assign _T_93 = sourceA_io_req_ready | _T_92; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100280.4]
  assign _T_94 = _T_91 & _T_93; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100281.4]
  assign _T_95 = ~abc_mshrs_1_io_schedule_bits_b_valid; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100282.4]
  assign _T_96 = sourceB_io_req_ready | _T_95; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100283.4]
  assign _T_97 = _T_94 & _T_96; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100284.4]
  assign _T_98 = ~abc_mshrs_1_io_schedule_bits_c_valid; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100285.4]
  assign _T_99 = sourceC_io_req_ready | _T_98; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100286.4]
  assign _T_100 = _T_97 & _T_99; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100287.4]
  assign _T_101 = ~abc_mshrs_1_io_schedule_bits_d_valid; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100288.4]
  assign _T_102 = sourceD_io_req_ready | _T_101; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100289.4]
  assign _T_103 = _T_100 & _T_102; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100290.4]
  assign _T_104 = ~abc_mshrs_1_io_schedule_bits_e_valid; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100291.4]
  assign _T_105 = sourceE_io_req_ready | _T_104; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100292.4]
  assign _T_106 = _T_103 & _T_105; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100293.4]
  assign _T_107 = ~abc_mshrs_1_io_schedule_bits_x_valid; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100294.4]
  assign _T_108 = sourceX_io_req_ready | _T_107; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100295.4]
  assign _T_109 = _T_106 & _T_108; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100296.4]
  assign _T_110 = ~abc_mshrs_1_io_schedule_bits_dir_valid; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100297.4]
  assign _T_111 = directory_io_write_ready | _T_110; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100298.4]
  assign _T_112 = _T_109 & _T_111; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100299.4]
  assign _T_113 = ~mshr_stall_2; // @[Scheduler.scala 105:28:chipyard.TestHarness.RocketConfig.fir@100300.4]
  assign _T_114 = abc_mshrs_2_io_schedule_valid & _T_113; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100301.4]
  assign _T_115 = ~abc_mshrs_2_io_schedule_bits_a_valid; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100302.4]
  assign _T_116 = sourceA_io_req_ready | _T_115; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100303.4]
  assign _T_117 = _T_114 & _T_116; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100304.4]
  assign _T_118 = ~abc_mshrs_2_io_schedule_bits_b_valid; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100305.4]
  assign _T_119 = sourceB_io_req_ready | _T_118; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100306.4]
  assign _T_120 = _T_117 & _T_119; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100307.4]
  assign _T_121 = ~abc_mshrs_2_io_schedule_bits_c_valid; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100308.4]
  assign _T_122 = sourceC_io_req_ready | _T_121; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100309.4]
  assign _T_123 = _T_120 & _T_122; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100310.4]
  assign _T_124 = ~abc_mshrs_2_io_schedule_bits_d_valid; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100311.4]
  assign _T_125 = sourceD_io_req_ready | _T_124; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100312.4]
  assign _T_126 = _T_123 & _T_125; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100313.4]
  assign _T_127 = ~abc_mshrs_2_io_schedule_bits_e_valid; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100314.4]
  assign _T_128 = sourceE_io_req_ready | _T_127; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100315.4]
  assign _T_129 = _T_126 & _T_128; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100316.4]
  assign _T_130 = ~abc_mshrs_2_io_schedule_bits_x_valid; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100317.4]
  assign _T_131 = sourceX_io_req_ready | _T_130; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100318.4]
  assign _T_132 = _T_129 & _T_131; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100319.4]
  assign _T_133 = ~abc_mshrs_2_io_schedule_bits_dir_valid; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100320.4]
  assign _T_134 = directory_io_write_ready | _T_133; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100321.4]
  assign _T_135 = _T_132 & _T_134; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100322.4]
  assign _T_136 = ~mshr_stall_3; // @[Scheduler.scala 105:28:chipyard.TestHarness.RocketConfig.fir@100323.4]
  assign _T_137 = abc_mshrs_3_io_schedule_valid & _T_136; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100324.4]
  assign _T_138 = ~abc_mshrs_3_io_schedule_bits_a_valid; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100325.4]
  assign _T_139 = sourceA_io_req_ready | _T_138; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100326.4]
  assign _T_140 = _T_137 & _T_139; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100327.4]
  assign _T_141 = ~abc_mshrs_3_io_schedule_bits_b_valid; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100328.4]
  assign _T_142 = sourceB_io_req_ready | _T_141; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100329.4]
  assign _T_143 = _T_140 & _T_142; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100330.4]
  assign _T_144 = ~abc_mshrs_3_io_schedule_bits_c_valid; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100331.4]
  assign _T_145 = sourceC_io_req_ready | _T_144; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100332.4]
  assign _T_146 = _T_143 & _T_145; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100333.4]
  assign _T_147 = ~abc_mshrs_3_io_schedule_bits_d_valid; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100334.4]
  assign _T_148 = sourceD_io_req_ready | _T_147; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100335.4]
  assign _T_149 = _T_146 & _T_148; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100336.4]
  assign _T_150 = ~abc_mshrs_3_io_schedule_bits_e_valid; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100337.4]
  assign _T_151 = sourceE_io_req_ready | _T_150; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100338.4]
  assign _T_152 = _T_149 & _T_151; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100339.4]
  assign _T_153 = ~abc_mshrs_3_io_schedule_bits_x_valid; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100340.4]
  assign _T_154 = sourceX_io_req_ready | _T_153; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100341.4]
  assign _T_155 = _T_152 & _T_154; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100342.4]
  assign _T_156 = ~abc_mshrs_3_io_schedule_bits_dir_valid; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100343.4]
  assign _T_157 = directory_io_write_ready | _T_156; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100344.4]
  assign _T_158 = _T_155 & _T_157; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100345.4]
  assign _T_159 = ~mshr_stall_4; // @[Scheduler.scala 105:28:chipyard.TestHarness.RocketConfig.fir@100346.4]
  assign _T_160 = abc_mshrs_4_io_schedule_valid & _T_159; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100347.4]
  assign _T_161 = ~abc_mshrs_4_io_schedule_bits_a_valid; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100348.4]
  assign _T_162 = sourceA_io_req_ready | _T_161; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100349.4]
  assign _T_163 = _T_160 & _T_162; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100350.4]
  assign _T_164 = ~abc_mshrs_4_io_schedule_bits_b_valid; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100351.4]
  assign _T_165 = sourceB_io_req_ready | _T_164; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100352.4]
  assign _T_166 = _T_163 & _T_165; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100353.4]
  assign _T_167 = ~abc_mshrs_4_io_schedule_bits_c_valid; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100354.4]
  assign _T_168 = sourceC_io_req_ready | _T_167; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100355.4]
  assign _T_169 = _T_166 & _T_168; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100356.4]
  assign _T_170 = ~abc_mshrs_4_io_schedule_bits_d_valid; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100357.4]
  assign _T_171 = sourceD_io_req_ready | _T_170; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100358.4]
  assign _T_172 = _T_169 & _T_171; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100359.4]
  assign _T_173 = ~abc_mshrs_4_io_schedule_bits_e_valid; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100360.4]
  assign _T_174 = sourceE_io_req_ready | _T_173; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100361.4]
  assign _T_175 = _T_172 & _T_174; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100362.4]
  assign _T_176 = ~abc_mshrs_4_io_schedule_bits_x_valid; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100363.4]
  assign _T_177 = sourceX_io_req_ready | _T_176; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100364.4]
  assign _T_178 = _T_175 & _T_177; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100365.4]
  assign _T_179 = ~abc_mshrs_4_io_schedule_bits_dir_valid; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100366.4]
  assign _T_180 = directory_io_write_ready | _T_179; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100367.4]
  assign _T_181 = _T_178 & _T_180; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100368.4]
  assign _T_182 = ~mshr_stall_5; // @[Scheduler.scala 105:28:chipyard.TestHarness.RocketConfig.fir@100369.4]
  assign _T_183 = bc_mshr_io_schedule_valid & _T_182; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100370.4]
  assign _T_184 = ~bc_mshr_io_schedule_bits_a_valid; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100371.4]
  assign _T_185 = sourceA_io_req_ready | _T_184; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100372.4]
  assign _T_186 = _T_183 & _T_185; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100373.4]
  assign _T_187 = ~bc_mshr_io_schedule_bits_b_valid; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100374.4]
  assign _T_188 = sourceB_io_req_ready | _T_187; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100375.4]
  assign _T_189 = _T_186 & _T_188; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100376.4]
  assign _T_190 = ~bc_mshr_io_schedule_bits_c_valid; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100377.4]
  assign _T_191 = sourceC_io_req_ready | _T_190; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100378.4]
  assign _T_192 = _T_189 & _T_191; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100379.4]
  assign _T_193 = ~bc_mshr_io_schedule_bits_d_valid; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100380.4]
  assign _T_194 = sourceD_io_req_ready | _T_193; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100381.4]
  assign _T_195 = _T_192 & _T_194; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100382.4]
  assign _T_196 = ~bc_mshr_io_schedule_bits_e_valid; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100383.4]
  assign _T_197 = sourceE_io_req_ready | _T_196; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100384.4]
  assign _T_198 = _T_195 & _T_197; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100385.4]
  assign _T_199 = ~bc_mshr_io_schedule_bits_x_valid; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100386.4]
  assign _T_200 = sourceX_io_req_ready | _T_199; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100387.4]
  assign _T_201 = _T_198 & _T_200; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100388.4]
  assign _T_202 = ~bc_mshr_io_schedule_bits_dir_valid; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100389.4]
  assign _T_203 = directory_io_write_ready | _T_202; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100390.4]
  assign _T_204 = _T_201 & _T_203; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100391.4]
  assign _T_206 = c_mshr_io_schedule_valid; // @[Scheduler.scala 105:25:chipyard.TestHarness.RocketConfig.fir@100393.4]
  assign _T_207 = ~c_mshr_io_schedule_bits_a_valid; // @[Scheduler.scala 106:32:chipyard.TestHarness.RocketConfig.fir@100394.4]
  assign _T_208 = sourceA_io_req_ready | _T_207; // @[Scheduler.scala 106:29:chipyard.TestHarness.RocketConfig.fir@100395.4]
  assign _T_209 = _T_206 & _T_208; // @[Scheduler.scala 105:31:chipyard.TestHarness.RocketConfig.fir@100396.4]
  assign _T_210 = ~c_mshr_io_schedule_bits_b_valid; // @[Scheduler.scala 107:32:chipyard.TestHarness.RocketConfig.fir@100397.4]
  assign _T_211 = sourceB_io_req_ready | _T_210; // @[Scheduler.scala 107:29:chipyard.TestHarness.RocketConfig.fir@100398.4]
  assign _T_212 = _T_209 & _T_211; // @[Scheduler.scala 106:61:chipyard.TestHarness.RocketConfig.fir@100399.4]
  assign _T_213 = ~c_mshr_io_schedule_bits_c_valid; // @[Scheduler.scala 108:32:chipyard.TestHarness.RocketConfig.fir@100400.4]
  assign _T_214 = sourceC_io_req_ready | _T_213; // @[Scheduler.scala 108:29:chipyard.TestHarness.RocketConfig.fir@100401.4]
  assign _T_215 = _T_212 & _T_214; // @[Scheduler.scala 107:61:chipyard.TestHarness.RocketConfig.fir@100402.4]
  assign _T_216 = ~c_mshr_io_schedule_bits_d_valid; // @[Scheduler.scala 109:32:chipyard.TestHarness.RocketConfig.fir@100403.4]
  assign _T_217 = sourceD_io_req_ready | _T_216; // @[Scheduler.scala 109:29:chipyard.TestHarness.RocketConfig.fir@100404.4]
  assign _T_218 = _T_215 & _T_217; // @[Scheduler.scala 108:61:chipyard.TestHarness.RocketConfig.fir@100405.4]
  assign _T_219 = ~c_mshr_io_schedule_bits_e_valid; // @[Scheduler.scala 110:32:chipyard.TestHarness.RocketConfig.fir@100406.4]
  assign _T_220 = sourceE_io_req_ready | _T_219; // @[Scheduler.scala 110:29:chipyard.TestHarness.RocketConfig.fir@100407.4]
  assign _T_221 = _T_218 & _T_220; // @[Scheduler.scala 109:61:chipyard.TestHarness.RocketConfig.fir@100408.4]
  assign _T_222 = ~c_mshr_io_schedule_bits_x_valid; // @[Scheduler.scala 111:32:chipyard.TestHarness.RocketConfig.fir@100409.4]
  assign _T_223 = sourceX_io_req_ready | _T_222; // @[Scheduler.scala 111:29:chipyard.TestHarness.RocketConfig.fir@100410.4]
  assign _T_224 = _T_221 & _T_223; // @[Scheduler.scala 110:61:chipyard.TestHarness.RocketConfig.fir@100411.4]
  assign _T_225 = ~c_mshr_io_schedule_bits_dir_valid; // @[Scheduler.scala 112:36:chipyard.TestHarness.RocketConfig.fir@100412.4]
  assign _T_226 = directory_io_write_ready | _T_225; // @[Scheduler.scala 112:33:chipyard.TestHarness.RocketConfig.fir@100413.4]
  assign _T_227 = _T_224 & _T_226; // @[Scheduler.scala 111:61:chipyard.TestHarness.RocketConfig.fir@100414.4]
  assign mshr_request = {_T_227,_T_204,_T_181,_T_158,_T_135,_T_112,_T_89}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@100420.4]
  assign _T_233 = mshr_request & robin_filter; // @[Scheduler.scala 117:54:chipyard.TestHarness.RocketConfig.fir@100422.4]
  assign robin_request = {_T_227,_T_204,_T_181,_T_158,_T_135,_T_112,_T_89,_T_233}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@100423.4]
  assign _T_234 = {robin_request, 1'h0}; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@100424.4]
  assign _T_236 = robin_request | _T_234[13:0]; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@100426.4]
  assign _T_237 = {_T_236, 2'h0}; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@100427.4]
  assign _T_239 = _T_236 | _T_237[13:0]; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@100429.4]
  assign _T_240 = {_T_239, 4'h0}; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@100430.4]
  assign _T_242 = _T_239 | _T_240[13:0]; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@100432.4]
  assign _T_243 = {_T_242, 8'h0}; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@100433.4]
  assign _T_245 = _T_242 | _T_243[13:0]; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@100435.4]
  assign _T_247 = {_T_245, 1'h0}; // @[Scheduler.scala 118:48:chipyard.TestHarness.RocketConfig.fir@100437.4]
  assign _T_248 = ~_T_247; // @[Scheduler.scala 118:24:chipyard.TestHarness.RocketConfig.fir@100438.4]
  assign _GEN_141 = {{1'd0}, robin_request}; // @[Scheduler.scala 118:54:chipyard.TestHarness.RocketConfig.fir@100439.4]
  assign mshr_selectOH2 = _T_248 & _GEN_141; // @[Scheduler.scala 118:54:chipyard.TestHarness.RocketConfig.fir@100439.4]
  assign mshr_selectOH = mshr_selectOH2[13:7] | mshr_selectOH2[6:0]; // @[Scheduler.scala 119:70:chipyard.TestHarness.RocketConfig.fir@100442.4]
  assign _T_253 = |mshr_selectOH[6:4]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@100445.4]
  assign _GEN_142 = {{1'd0}, mshr_selectOH[6:4]}; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@100446.4]
  assign _T_254 = _GEN_142 | mshr_selectOH[3:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@100446.4]
  assign _T_257 = |_T_254[3:2]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@100449.4]
  assign _T_258 = _T_254[3:2] | _T_254[1:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@100450.4]
  assign _T_260 = {_T_257,_T_258[1]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@100452.4]
  assign mshr_select = {_T_253,_T_257,_T_258[1]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@100453.4]
  assign _T_271 = {abc_mshrs_0_io_schedule_bits_dir_bits_data_dirty,abc_mshrs_0_io_schedule_bits_dir_bits_data_state,abc_mshrs_0_io_schedule_bits_dir_bits_data_clients,abc_mshrs_0_io_schedule_bits_dir_bits_data_tag,abc_mshrs_0_io_schedule_bits_reload}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100464.4]
  assign _T_277 = {abc_mshrs_0_io_schedule_bits_e_bits_sink,abc_mshrs_0_io_schedule_bits_x_valid,1'h0,abc_mshrs_0_io_schedule_bits_dir_valid,abc_mshrs_0_io_schedule_bits_dir_bits_set,abc_mshrs_0_io_schedule_bits_dir_bits_way,_T_271}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100470.4]
  assign _T_282 = {abc_mshrs_0_io_schedule_bits_d_bits_put,abc_mshrs_0_io_schedule_bits_d_bits_set,3'h0,abc_mshrs_0_io_schedule_bits_d_bits_way,abc_mshrs_0_io_schedule_bits_d_bits_bad,abc_mshrs_0_io_schedule_bits_e_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100475.4]
  assign _T_289 = {abc_mshrs_0_io_schedule_bits_d_bits_opcode,abc_mshrs_0_io_schedule_bits_d_bits_param,abc_mshrs_0_io_schedule_bits_d_bits_size,abc_mshrs_0_io_schedule_bits_d_bits_source,abc_mshrs_0_io_schedule_bits_d_bits_tag,abc_mshrs_0_io_schedule_bits_d_bits_offset,_T_282,_T_277}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100482.4]
  assign _T_294 = {abc_mshrs_0_io_schedule_bits_c_bits_dirty,abc_mshrs_0_io_schedule_bits_d_valid,abc_mshrs_0_io_schedule_bits_d_bits_prio_2,abc_mshrs_0_io_schedule_bits_d_bits_prio_1,abc_mshrs_0_io_schedule_bits_d_bits_prio_0,abc_mshrs_0_io_schedule_bits_d_bits_control}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100487.4]
  assign _T_300 = {abc_mshrs_0_io_schedule_bits_c_bits_opcode,abc_mshrs_0_io_schedule_bits_c_bits_param,3'h0,abc_mshrs_0_io_schedule_bits_c_bits_tag,abc_mshrs_0_io_schedule_bits_c_bits_set,abc_mshrs_0_io_schedule_bits_c_bits_way,_T_294}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100493.4]
  assign _T_305 = {abc_mshrs_0_io_schedule_bits_b_valid,abc_mshrs_0_io_schedule_bits_b_bits_param,abc_mshrs_0_io_schedule_bits_b_bits_tag,abc_mshrs_0_io_schedule_bits_b_bits_set,abc_mshrs_0_io_schedule_bits_b_bits_clients,abc_mshrs_0_io_schedule_bits_c_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100498.4]
  assign _T_313 = {abc_mshrs_0_io_schedule_bits_a_valid,abc_mshrs_0_io_schedule_bits_a_bits_tag,abc_mshrs_0_io_schedule_bits_a_bits_set,abc_mshrs_0_io_schedule_bits_a_bits_param,3'h0,abc_mshrs_0_io_schedule_bits_a_bits_block,_T_305,_T_300,_T_289}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100506.4]
  assign _T_314 = mshr_selectOH[0] ? _T_313 : 188'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100507.4]
  assign _T_318 = {abc_mshrs_1_io_schedule_bits_dir_bits_data_dirty,abc_mshrs_1_io_schedule_bits_dir_bits_data_state,abc_mshrs_1_io_schedule_bits_dir_bits_data_clients,abc_mshrs_1_io_schedule_bits_dir_bits_data_tag,abc_mshrs_1_io_schedule_bits_reload}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100511.4]
  assign _T_324 = {abc_mshrs_1_io_schedule_bits_e_bits_sink,abc_mshrs_1_io_schedule_bits_x_valid,1'h0,abc_mshrs_1_io_schedule_bits_dir_valid,abc_mshrs_1_io_schedule_bits_dir_bits_set,abc_mshrs_1_io_schedule_bits_dir_bits_way,_T_318}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100517.4]
  assign _T_329 = {abc_mshrs_1_io_schedule_bits_d_bits_put,abc_mshrs_1_io_schedule_bits_d_bits_set,3'h0,abc_mshrs_1_io_schedule_bits_d_bits_way,abc_mshrs_1_io_schedule_bits_d_bits_bad,abc_mshrs_1_io_schedule_bits_e_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100522.4]
  assign _T_336 = {abc_mshrs_1_io_schedule_bits_d_bits_opcode,abc_mshrs_1_io_schedule_bits_d_bits_param,abc_mshrs_1_io_schedule_bits_d_bits_size,abc_mshrs_1_io_schedule_bits_d_bits_source,abc_mshrs_1_io_schedule_bits_d_bits_tag,abc_mshrs_1_io_schedule_bits_d_bits_offset,_T_329,_T_324}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100529.4]
  assign _T_341 = {abc_mshrs_1_io_schedule_bits_c_bits_dirty,abc_mshrs_1_io_schedule_bits_d_valid,abc_mshrs_1_io_schedule_bits_d_bits_prio_2,abc_mshrs_1_io_schedule_bits_d_bits_prio_1,abc_mshrs_1_io_schedule_bits_d_bits_prio_0,abc_mshrs_1_io_schedule_bits_d_bits_control}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100534.4]
  assign _T_347 = {abc_mshrs_1_io_schedule_bits_c_bits_opcode,abc_mshrs_1_io_schedule_bits_c_bits_param,3'h0,abc_mshrs_1_io_schedule_bits_c_bits_tag,abc_mshrs_1_io_schedule_bits_c_bits_set,abc_mshrs_1_io_schedule_bits_c_bits_way,_T_341}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100540.4]
  assign _T_352 = {abc_mshrs_1_io_schedule_bits_b_valid,abc_mshrs_1_io_schedule_bits_b_bits_param,abc_mshrs_1_io_schedule_bits_b_bits_tag,abc_mshrs_1_io_schedule_bits_b_bits_set,abc_mshrs_1_io_schedule_bits_b_bits_clients,abc_mshrs_1_io_schedule_bits_c_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100545.4]
  assign _T_360 = {abc_mshrs_1_io_schedule_bits_a_valid,abc_mshrs_1_io_schedule_bits_a_bits_tag,abc_mshrs_1_io_schedule_bits_a_bits_set,abc_mshrs_1_io_schedule_bits_a_bits_param,3'h0,abc_mshrs_1_io_schedule_bits_a_bits_block,_T_352,_T_347,_T_336}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100553.4]
  assign _T_361 = mshr_selectOH[1] ? _T_360 : 188'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100554.4]
  assign _T_365 = {abc_mshrs_2_io_schedule_bits_dir_bits_data_dirty,abc_mshrs_2_io_schedule_bits_dir_bits_data_state,abc_mshrs_2_io_schedule_bits_dir_bits_data_clients,abc_mshrs_2_io_schedule_bits_dir_bits_data_tag,abc_mshrs_2_io_schedule_bits_reload}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100558.4]
  assign _T_371 = {abc_mshrs_2_io_schedule_bits_e_bits_sink,abc_mshrs_2_io_schedule_bits_x_valid,1'h0,abc_mshrs_2_io_schedule_bits_dir_valid,abc_mshrs_2_io_schedule_bits_dir_bits_set,abc_mshrs_2_io_schedule_bits_dir_bits_way,_T_365}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100564.4]
  assign _T_376 = {abc_mshrs_2_io_schedule_bits_d_bits_put,abc_mshrs_2_io_schedule_bits_d_bits_set,3'h0,abc_mshrs_2_io_schedule_bits_d_bits_way,abc_mshrs_2_io_schedule_bits_d_bits_bad,abc_mshrs_2_io_schedule_bits_e_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100569.4]
  assign _T_383 = {abc_mshrs_2_io_schedule_bits_d_bits_opcode,abc_mshrs_2_io_schedule_bits_d_bits_param,abc_mshrs_2_io_schedule_bits_d_bits_size,abc_mshrs_2_io_schedule_bits_d_bits_source,abc_mshrs_2_io_schedule_bits_d_bits_tag,abc_mshrs_2_io_schedule_bits_d_bits_offset,_T_376,_T_371}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100576.4]
  assign _T_388 = {abc_mshrs_2_io_schedule_bits_c_bits_dirty,abc_mshrs_2_io_schedule_bits_d_valid,abc_mshrs_2_io_schedule_bits_d_bits_prio_2,abc_mshrs_2_io_schedule_bits_d_bits_prio_1,abc_mshrs_2_io_schedule_bits_d_bits_prio_0,abc_mshrs_2_io_schedule_bits_d_bits_control}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100581.4]
  assign _T_394 = {abc_mshrs_2_io_schedule_bits_c_bits_opcode,abc_mshrs_2_io_schedule_bits_c_bits_param,3'h0,abc_mshrs_2_io_schedule_bits_c_bits_tag,abc_mshrs_2_io_schedule_bits_c_bits_set,abc_mshrs_2_io_schedule_bits_c_bits_way,_T_388}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100587.4]
  assign _T_399 = {abc_mshrs_2_io_schedule_bits_b_valid,abc_mshrs_2_io_schedule_bits_b_bits_param,abc_mshrs_2_io_schedule_bits_b_bits_tag,abc_mshrs_2_io_schedule_bits_b_bits_set,abc_mshrs_2_io_schedule_bits_b_bits_clients,abc_mshrs_2_io_schedule_bits_c_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100592.4]
  assign _T_407 = {abc_mshrs_2_io_schedule_bits_a_valid,abc_mshrs_2_io_schedule_bits_a_bits_tag,abc_mshrs_2_io_schedule_bits_a_bits_set,abc_mshrs_2_io_schedule_bits_a_bits_param,3'h0,abc_mshrs_2_io_schedule_bits_a_bits_block,_T_399,_T_394,_T_383}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100600.4]
  assign _T_408 = mshr_selectOH[2] ? _T_407 : 188'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100601.4]
  assign _T_412 = {abc_mshrs_3_io_schedule_bits_dir_bits_data_dirty,abc_mshrs_3_io_schedule_bits_dir_bits_data_state,abc_mshrs_3_io_schedule_bits_dir_bits_data_clients,abc_mshrs_3_io_schedule_bits_dir_bits_data_tag,abc_mshrs_3_io_schedule_bits_reload}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100605.4]
  assign _T_418 = {abc_mshrs_3_io_schedule_bits_e_bits_sink,abc_mshrs_3_io_schedule_bits_x_valid,1'h0,abc_mshrs_3_io_schedule_bits_dir_valid,abc_mshrs_3_io_schedule_bits_dir_bits_set,abc_mshrs_3_io_schedule_bits_dir_bits_way,_T_412}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100611.4]
  assign _T_423 = {abc_mshrs_3_io_schedule_bits_d_bits_put,abc_mshrs_3_io_schedule_bits_d_bits_set,3'h0,abc_mshrs_3_io_schedule_bits_d_bits_way,abc_mshrs_3_io_schedule_bits_d_bits_bad,abc_mshrs_3_io_schedule_bits_e_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100616.4]
  assign _T_430 = {abc_mshrs_3_io_schedule_bits_d_bits_opcode,abc_mshrs_3_io_schedule_bits_d_bits_param,abc_mshrs_3_io_schedule_bits_d_bits_size,abc_mshrs_3_io_schedule_bits_d_bits_source,abc_mshrs_3_io_schedule_bits_d_bits_tag,abc_mshrs_3_io_schedule_bits_d_bits_offset,_T_423,_T_418}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100623.4]
  assign _T_435 = {abc_mshrs_3_io_schedule_bits_c_bits_dirty,abc_mshrs_3_io_schedule_bits_d_valid,abc_mshrs_3_io_schedule_bits_d_bits_prio_2,abc_mshrs_3_io_schedule_bits_d_bits_prio_1,abc_mshrs_3_io_schedule_bits_d_bits_prio_0,abc_mshrs_3_io_schedule_bits_d_bits_control}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100628.4]
  assign _T_441 = {abc_mshrs_3_io_schedule_bits_c_bits_opcode,abc_mshrs_3_io_schedule_bits_c_bits_param,3'h0,abc_mshrs_3_io_schedule_bits_c_bits_tag,abc_mshrs_3_io_schedule_bits_c_bits_set,abc_mshrs_3_io_schedule_bits_c_bits_way,_T_435}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100634.4]
  assign _T_446 = {abc_mshrs_3_io_schedule_bits_b_valid,abc_mshrs_3_io_schedule_bits_b_bits_param,abc_mshrs_3_io_schedule_bits_b_bits_tag,abc_mshrs_3_io_schedule_bits_b_bits_set,abc_mshrs_3_io_schedule_bits_b_bits_clients,abc_mshrs_3_io_schedule_bits_c_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100639.4]
  assign _T_454 = {abc_mshrs_3_io_schedule_bits_a_valid,abc_mshrs_3_io_schedule_bits_a_bits_tag,abc_mshrs_3_io_schedule_bits_a_bits_set,abc_mshrs_3_io_schedule_bits_a_bits_param,3'h0,abc_mshrs_3_io_schedule_bits_a_bits_block,_T_446,_T_441,_T_430}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100647.4]
  assign _T_455 = mshr_selectOH[3] ? _T_454 : 188'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100648.4]
  assign _T_459 = {abc_mshrs_4_io_schedule_bits_dir_bits_data_dirty,abc_mshrs_4_io_schedule_bits_dir_bits_data_state,abc_mshrs_4_io_schedule_bits_dir_bits_data_clients,abc_mshrs_4_io_schedule_bits_dir_bits_data_tag,abc_mshrs_4_io_schedule_bits_reload}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100652.4]
  assign _T_465 = {abc_mshrs_4_io_schedule_bits_e_bits_sink,abc_mshrs_4_io_schedule_bits_x_valid,1'h0,abc_mshrs_4_io_schedule_bits_dir_valid,abc_mshrs_4_io_schedule_bits_dir_bits_set,abc_mshrs_4_io_schedule_bits_dir_bits_way,_T_459}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100658.4]
  assign _T_470 = {abc_mshrs_4_io_schedule_bits_d_bits_put,abc_mshrs_4_io_schedule_bits_d_bits_set,3'h0,abc_mshrs_4_io_schedule_bits_d_bits_way,abc_mshrs_4_io_schedule_bits_d_bits_bad,abc_mshrs_4_io_schedule_bits_e_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100663.4]
  assign _T_477 = {abc_mshrs_4_io_schedule_bits_d_bits_opcode,abc_mshrs_4_io_schedule_bits_d_bits_param,abc_mshrs_4_io_schedule_bits_d_bits_size,abc_mshrs_4_io_schedule_bits_d_bits_source,abc_mshrs_4_io_schedule_bits_d_bits_tag,abc_mshrs_4_io_schedule_bits_d_bits_offset,_T_470,_T_465}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100670.4]
  assign _T_482 = {abc_mshrs_4_io_schedule_bits_c_bits_dirty,abc_mshrs_4_io_schedule_bits_d_valid,abc_mshrs_4_io_schedule_bits_d_bits_prio_2,abc_mshrs_4_io_schedule_bits_d_bits_prio_1,abc_mshrs_4_io_schedule_bits_d_bits_prio_0,abc_mshrs_4_io_schedule_bits_d_bits_control}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100675.4]
  assign _T_488 = {abc_mshrs_4_io_schedule_bits_c_bits_opcode,abc_mshrs_4_io_schedule_bits_c_bits_param,3'h0,abc_mshrs_4_io_schedule_bits_c_bits_tag,abc_mshrs_4_io_schedule_bits_c_bits_set,abc_mshrs_4_io_schedule_bits_c_bits_way,_T_482}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100681.4]
  assign _T_493 = {abc_mshrs_4_io_schedule_bits_b_valid,abc_mshrs_4_io_schedule_bits_b_bits_param,abc_mshrs_4_io_schedule_bits_b_bits_tag,abc_mshrs_4_io_schedule_bits_b_bits_set,abc_mshrs_4_io_schedule_bits_b_bits_clients,abc_mshrs_4_io_schedule_bits_c_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100686.4]
  assign _T_501 = {abc_mshrs_4_io_schedule_bits_a_valid,abc_mshrs_4_io_schedule_bits_a_bits_tag,abc_mshrs_4_io_schedule_bits_a_bits_set,abc_mshrs_4_io_schedule_bits_a_bits_param,3'h0,abc_mshrs_4_io_schedule_bits_a_bits_block,_T_493,_T_488,_T_477}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100694.4]
  assign _T_502 = mshr_selectOH[4] ? _T_501 : 188'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100695.4]
  assign _T_506 = {bc_mshr_io_schedule_bits_dir_bits_data_dirty,bc_mshr_io_schedule_bits_dir_bits_data_state,bc_mshr_io_schedule_bits_dir_bits_data_clients,bc_mshr_io_schedule_bits_dir_bits_data_tag,bc_mshr_io_schedule_bits_reload}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100699.4]
  assign _T_512 = {bc_mshr_io_schedule_bits_e_bits_sink,bc_mshr_io_schedule_bits_x_valid,1'h0,bc_mshr_io_schedule_bits_dir_valid,bc_mshr_io_schedule_bits_dir_bits_set,bc_mshr_io_schedule_bits_dir_bits_way,_T_506}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100705.4]
  assign _T_517 = {bc_mshr_io_schedule_bits_d_bits_put,bc_mshr_io_schedule_bits_d_bits_set,3'h0,bc_mshr_io_schedule_bits_d_bits_way,bc_mshr_io_schedule_bits_d_bits_bad,bc_mshr_io_schedule_bits_e_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100710.4]
  assign _T_524 = {bc_mshr_io_schedule_bits_d_bits_opcode,bc_mshr_io_schedule_bits_d_bits_param,bc_mshr_io_schedule_bits_d_bits_size,bc_mshr_io_schedule_bits_d_bits_source,bc_mshr_io_schedule_bits_d_bits_tag,bc_mshr_io_schedule_bits_d_bits_offset,_T_517,_T_512}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100717.4]
  assign _T_529 = {bc_mshr_io_schedule_bits_c_bits_dirty,bc_mshr_io_schedule_bits_d_valid,bc_mshr_io_schedule_bits_d_bits_prio_2,bc_mshr_io_schedule_bits_d_bits_prio_1,bc_mshr_io_schedule_bits_d_bits_prio_0,bc_mshr_io_schedule_bits_d_bits_control}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100722.4]
  assign _T_535 = {bc_mshr_io_schedule_bits_c_bits_opcode,bc_mshr_io_schedule_bits_c_bits_param,3'h0,bc_mshr_io_schedule_bits_c_bits_tag,bc_mshr_io_schedule_bits_c_bits_set,bc_mshr_io_schedule_bits_c_bits_way,_T_529}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100728.4]
  assign _T_540 = {bc_mshr_io_schedule_bits_b_valid,bc_mshr_io_schedule_bits_b_bits_param,bc_mshr_io_schedule_bits_b_bits_tag,bc_mshr_io_schedule_bits_b_bits_set,bc_mshr_io_schedule_bits_b_bits_clients,bc_mshr_io_schedule_bits_c_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100733.4]
  assign _T_548 = {bc_mshr_io_schedule_bits_a_valid,bc_mshr_io_schedule_bits_a_bits_tag,bc_mshr_io_schedule_bits_a_bits_set,bc_mshr_io_schedule_bits_a_bits_param,3'h0,bc_mshr_io_schedule_bits_a_bits_block,_T_540,_T_535,_T_524}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100741.4]
  assign _T_549 = mshr_selectOH[5] ? _T_548 : 188'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100742.4]
  assign _T_553 = {c_mshr_io_schedule_bits_dir_bits_data_dirty,c_mshr_io_schedule_bits_dir_bits_data_state,c_mshr_io_schedule_bits_dir_bits_data_clients,c_mshr_io_schedule_bits_dir_bits_data_tag,c_mshr_io_schedule_bits_reload}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100746.4]
  assign _T_559 = {c_mshr_io_schedule_bits_e_bits_sink,c_mshr_io_schedule_bits_x_valid,1'h0,c_mshr_io_schedule_bits_dir_valid,c_mshr_io_schedule_bits_dir_bits_set,c_mshr_io_schedule_bits_dir_bits_way,_T_553}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100752.4]
  assign _T_564 = {c_mshr_io_schedule_bits_d_bits_put,c_mshr_io_schedule_bits_d_bits_set,3'h0,c_mshr_io_schedule_bits_d_bits_way,c_mshr_io_schedule_bits_d_bits_bad,c_mshr_io_schedule_bits_e_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100757.4]
  assign _T_571 = {c_mshr_io_schedule_bits_d_bits_opcode,c_mshr_io_schedule_bits_d_bits_param,c_mshr_io_schedule_bits_d_bits_size,c_mshr_io_schedule_bits_d_bits_source,c_mshr_io_schedule_bits_d_bits_tag,c_mshr_io_schedule_bits_d_bits_offset,_T_564,_T_559}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100764.4]
  assign _T_576 = {c_mshr_io_schedule_bits_c_bits_dirty,c_mshr_io_schedule_bits_d_valid,c_mshr_io_schedule_bits_d_bits_prio_2,c_mshr_io_schedule_bits_d_bits_prio_1,c_mshr_io_schedule_bits_d_bits_prio_0,c_mshr_io_schedule_bits_d_bits_control}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100769.4]
  assign _T_582 = {c_mshr_io_schedule_bits_c_bits_opcode,c_mshr_io_schedule_bits_c_bits_param,3'h0,c_mshr_io_schedule_bits_c_bits_tag,c_mshr_io_schedule_bits_c_bits_set,c_mshr_io_schedule_bits_c_bits_way,_T_576}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100775.4]
  assign _T_587 = {c_mshr_io_schedule_bits_b_valid,c_mshr_io_schedule_bits_b_bits_param,c_mshr_io_schedule_bits_b_bits_tag,c_mshr_io_schedule_bits_b_bits_set,c_mshr_io_schedule_bits_b_bits_clients,c_mshr_io_schedule_bits_c_valid}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100780.4]
  assign _T_595 = {c_mshr_io_schedule_bits_a_valid,c_mshr_io_schedule_bits_a_bits_tag,c_mshr_io_schedule_bits_a_bits_set,c_mshr_io_schedule_bits_a_bits_param,3'h0,c_mshr_io_schedule_bits_a_bits_block,_T_587,_T_582,_T_571}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100788.4]
  assign _T_596 = mshr_selectOH[6] ? _T_595 : 188'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100789.4]
  assign _T_597 = _T_314 | _T_361; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100790.4]
  assign _T_598 = _T_597 | _T_408; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100791.4]
  assign _T_599 = _T_598 | _T_455; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100792.4]
  assign _T_600 = _T_599 | _T_502; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100793.4]
  assign _T_601 = _T_600 | _T_549; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100794.4]
  assign _T_602 = _T_601 | _T_596; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100795.4]
  assign schedule_reload = _T_602[0]; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100799.4]
  assign schedule_c_bits_opcode = _T_602[129:127]; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100867.4]
  assign _T_658 = mshr_selectOH[0] ? abc_mshrs_0_io_status_bits_tag : 12'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100900.4]
  assign _T_659 = mshr_selectOH[1] ? abc_mshrs_1_io_status_bits_tag : 12'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100901.4]
  assign _T_660 = mshr_selectOH[2] ? abc_mshrs_2_io_status_bits_tag : 12'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100902.4]
  assign _T_661 = mshr_selectOH[3] ? abc_mshrs_3_io_status_bits_tag : 12'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100903.4]
  assign _T_662 = mshr_selectOH[4] ? abc_mshrs_4_io_status_bits_tag : 12'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100904.4]
  assign _T_663 = mshr_selectOH[5] ? bc_mshr_io_status_bits_tag : 12'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100905.4]
  assign _T_664 = mshr_selectOH[6] ? c_mshr_io_status_bits_tag : 12'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100906.4]
  assign _T_665 = _T_658 | _T_659; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100907.4]
  assign _T_666 = _T_665 | _T_660; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100908.4]
  assign _T_667 = _T_666 | _T_661; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100909.4]
  assign _T_668 = _T_667 | _T_662; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100910.4]
  assign _T_669 = _T_668 | _T_663; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100911.4]
  assign scheduleTag = _T_669 | _T_664; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100912.4]
  assign _T_678 = mshr_selectOH[0] ? abc_mshrs_0_io_status_bits_set : 10'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100922.4]
  assign _T_679 = mshr_selectOH[1] ? abc_mshrs_1_io_status_bits_set : 10'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100923.4]
  assign _T_680 = mshr_selectOH[2] ? abc_mshrs_2_io_status_bits_set : 10'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100924.4]
  assign _T_681 = mshr_selectOH[3] ? abc_mshrs_3_io_status_bits_set : 10'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100925.4]
  assign _T_682 = mshr_selectOH[4] ? abc_mshrs_4_io_status_bits_set : 10'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100926.4]
  assign _T_683 = mshr_selectOH[5] ? bc_mshr_io_status_bits_set : 10'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100927.4]
  assign _T_684 = mshr_selectOH[6] ? c_mshr_io_status_bits_set : 10'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100928.4]
  assign _T_685 = _T_678 | _T_679; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100929.4]
  assign _T_686 = _T_685 | _T_680; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100930.4]
  assign _T_687 = _T_686 | _T_681; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100931.4]
  assign _T_688 = _T_687 | _T_682; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100932.4]
  assign _T_689 = _T_688 | _T_683; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100933.4]
  assign scheduleSet = _T_689 | _T_684; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@100934.4]
  assign _T_691 = |mshr_request; // @[Scheduler.scala 126:25:chipyard.TestHarness.RocketConfig.fir@100937.4]
  assign _GEN_143 = {{1'd0}, mshr_selectOH[6:1]}; // @[package.scala 208:43:chipyard.TestHarness.RocketConfig.fir@100940.6]
  assign _T_693 = mshr_selectOH | _GEN_143; // @[package.scala 208:43:chipyard.TestHarness.RocketConfig.fir@100940.6]
  assign _GEN_144 = {{2'd0}, _T_693[6:2]}; // @[package.scala 208:43:chipyard.TestHarness.RocketConfig.fir@100942.6]
  assign _T_695 = _T_693 | _GEN_144; // @[package.scala 208:43:chipyard.TestHarness.RocketConfig.fir@100942.6]
  assign _GEN_145 = {{4'd0}, _T_695[6:4]}; // @[package.scala 208:43:chipyard.TestHarness.RocketConfig.fir@100944.6]
  assign _T_697 = _T_695 | _GEN_145; // @[package.scala 208:43:chipyard.TestHarness.RocketConfig.fir@100944.6]
  assign _T_699 = ~_T_697; // @[Scheduler.scala 126:47:chipyard.TestHarness.RocketConfig.fir@100946.6]
  assign _T_704 = mshr_selectOH[5] & bc_mshr_io_schedule_bits_dir_valid; // @[Scheduler.scala 146:37:chipyard.TestHarness.RocketConfig.fir@100967.4]
  assign _T_705 = bc_mshr_io_schedule_bits_dir_bits_data_state == 2'h0; // @[Scheduler.scala 146:123:chipyard.TestHarness.RocketConfig.fir@100968.4]
  assign _T_708 = bc_mshr_io_schedule_bits_dir_bits_data_state == 2'h1; // @[Scheduler.scala 147:123:chipyard.TestHarness.RocketConfig.fir@100972.4]
  assign _T_711 = mshr_selectOH[6] & c_mshr_io_schedule_bits_dir_valid; // @[Scheduler.scala 149:37:chipyard.TestHarness.RocketConfig.fir@100977.4]
  assign _T_713 = sinkA_io_req_valid | sinkX_io_req_valid; // @[Scheduler.scala 153:62:chipyard.TestHarness.RocketConfig.fir@100982.4]
  assign _T_714 = _T_713 | sinkC_io_req_valid; // @[Scheduler.scala 153:84:chipyard.TestHarness.RocketConfig.fir@100983.4]
  assign request_valid = directory_io_ready & _T_714; // @[Scheduler.scala 153:39:chipyard.TestHarness.RocketConfig.fir@100984.4]
  assign _T_716_control = sinkX_io_req_valid; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  assign _T_716_opcode = sinkX_io_req_valid ? 3'h0 : sinkA_io_req_bits_opcode; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  assign _T_716_param = sinkX_io_req_valid ? 3'h0 : sinkA_io_req_bits_param; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  assign _T_716_size = sinkX_io_req_valid ? 3'h6 : sinkA_io_req_bits_size; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  assign _T_716_source = sinkX_io_req_valid ? 3'h0 : sinkA_io_req_bits_source; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  assign _T_716_tag = sinkX_io_req_valid ? sinkX_io_req_bits_tag : sinkA_io_req_bits_tag; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  assign _T_716_offset = sinkX_io_req_valid ? 6'h0 : sinkA_io_req_bits_offset; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  assign _T_716_put = sinkX_io_req_valid ? 6'h0 : sinkA_io_req_bits_put; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  assign _T_716_set = sinkX_io_req_valid ? sinkX_io_req_bits_set : sinkA_io_req_bits_set; // @[Scheduler.scala 155:22:chipyard.TestHarness.RocketConfig.fir@100986.4]
  assign request_bits_prio_0 = sinkC_io_req_valid ? 1'h0 : 1'h1; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  assign request_bits_prio_2 = sinkC_io_req_valid; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  assign request_bits_control = sinkC_io_req_valid ? 1'h0 : _T_716_control; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  assign request_bits_opcode = sinkC_io_req_valid ? sinkC_io_req_bits_opcode : _T_716_opcode; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  assign request_bits_param = sinkC_io_req_valid ? sinkC_io_req_bits_param : _T_716_param; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  assign request_bits_size = sinkC_io_req_valid ? sinkC_io_req_bits_size : _T_716_size; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  assign request_bits_source = sinkC_io_req_valid ? sinkC_io_req_bits_source : _T_716_source; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  assign request_bits_tag = sinkC_io_req_valid ? sinkC_io_req_bits_tag : _T_716_tag; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  assign request_bits_offset = sinkC_io_req_valid ? sinkC_io_req_bits_offset : _T_716_offset; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  assign request_bits_put = sinkC_io_req_valid ? sinkC_io_req_bits_put : _T_716_put; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  assign request_bits_set = sinkC_io_req_valid ? sinkC_io_req_bits_set : _T_716_set; // @[Scheduler.scala 154:22:chipyard.TestHarness.RocketConfig.fir@100987.4]
  assign _T_739 = c_mshr_io_status_bits_set == request_bits_set; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101013.4]
  assign _T_740 = c_mshr_io_status_valid & _T_739; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101014.4]
  assign _T_737 = bc_mshr_io_status_bits_set == request_bits_set; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101011.4]
  assign _T_738 = bc_mshr_io_status_valid & _T_737; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101012.4]
  assign _T_735 = abc_mshrs_4_io_status_bits_set == request_bits_set; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101009.4]
  assign _T_736 = abc_mshrs_4_io_status_valid & _T_735; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101010.4]
  assign _T_733 = abc_mshrs_3_io_status_bits_set == request_bits_set; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101007.4]
  assign _T_734 = abc_mshrs_3_io_status_valid & _T_733; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101008.4]
  assign _T_731 = abc_mshrs_2_io_status_bits_set == request_bits_set; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101005.4]
  assign _T_732 = abc_mshrs_2_io_status_valid & _T_731; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101006.4]
  assign _T_729 = abc_mshrs_1_io_status_bits_set == request_bits_set; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101003.4]
  assign _T_730 = abc_mshrs_1_io_status_valid & _T_729; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101004.4]
  assign _T_727 = abc_mshrs_0_io_status_bits_set == request_bits_set; // @[Scheduler.scala 161:83:chipyard.TestHarness.RocketConfig.fir@101001.4]
  assign _T_728 = abc_mshrs_0_io_status_valid & _T_727; // @[Scheduler.scala 161:59:chipyard.TestHarness.RocketConfig.fir@101002.4]
  assign setMatches = {_T_740,_T_738,_T_736,_T_734,_T_732,_T_730,_T_728}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101020.4]
  assign _T_746 = |setMatches; // @[Scheduler.scala 162:30:chipyard.TestHarness.RocketConfig.fir@101021.4]
  assign alloc = ~_T_746; // @[Scheduler.scala 162:15:chipyard.TestHarness.RocketConfig.fir@101022.4]
  assign _T_849 = {mshr_selectOH,mshr_selectOH,mshr_selectOH}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101137.4]
  assign selected_requests = _T_849 & requests_io_valid; // @[Scheduler.scala 195:76:chipyard.TestHarness.RocketConfig.fir@101138.4]
  assign a_pop = |selected_requests[6:0]; // @[Scheduler.scala 196:82:chipyard.TestHarness.RocketConfig.fir@101140.4]
  assign b_pop = |selected_requests[13:7]; // @[Scheduler.scala 197:82:chipyard.TestHarness.RocketConfig.fir@101142.4]
  assign _T_862 = a_pop | b_pop; // @[Scheduler.scala 201:23:chipyard.TestHarness.RocketConfig.fir@101155.4]
  assign c_pop = |selected_requests[20:14]; // @[Scheduler.scala 198:82:chipyard.TestHarness.RocketConfig.fir@101144.4]
  assign may_pop = _T_862 | c_pop; // @[Scheduler.scala 201:32:chipyard.TestHarness.RocketConfig.fir@101156.4]
  assign _T_1062 = schedule_reload & may_pop; // @[Scheduler.scala 236:64:chipyard.TestHarness.RocketConfig.fir@101413.4]
  assign lb_tag_mismatch = scheduleTag != requests_io_data_tag; // @[Scheduler.scala 235:37:chipyard.TestHarness.RocketConfig.fir@101412.4]
  assign mshr_uses_directory_assuming_no_bypass = _T_1062 & lb_tag_mismatch; // @[Scheduler.scala 236:75:chipyard.TestHarness.RocketConfig.fir@101414.4]
  assign _T_1072 = ~mshr_uses_directory_assuming_no_bypass; // @[Scheduler.scala 247:16:chipyard.TestHarness.RocketConfig.fir@101429.4]
  assign _T_1073 = alloc & _T_1072; // @[Scheduler.scala 247:13:chipyard.TestHarness.RocketConfig.fir@101430.4]
  assign mshr_validOH = {c_mshr_io_status_valid,bc_mshr_io_status_valid,abc_mshrs_4_io_status_valid,abc_mshrs_3_io_status_valid,abc_mshrs_2_io_status_valid,abc_mshrs_1_io_status_valid,abc_mshrs_0_io_status_valid}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101424.4]
  assign _T_1070 = ~mshr_validOH; // @[Scheduler.scala 242:20:chipyard.TestHarness.RocketConfig.fir@101425.4]
  assign _T_831 = ~request_bits_prio_0; // @[Scheduler.scala 171:46:chipyard.TestHarness.RocketConfig.fir@101115.4]
  assign prioFilter = {request_bits_prio_2,_T_831,5'h1f}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101118.4]
  assign _T_1071 = _T_1070 & prioFilter; // @[Scheduler.scala 242:34:chipyard.TestHarness.RocketConfig.fir@101426.4]
  assign mshr_free = |_T_1071; // @[Scheduler.scala 242:51:chipyard.TestHarness.RocketConfig.fir@101427.4]
  assign _T_1074 = _T_1073 & mshr_free; // @[Scheduler.scala 247:56:chipyard.TestHarness.RocketConfig.fir@101431.4]
  assign _T_1079 = ~c_mshr_io_status_valid; // @[Scheduler.scala 248:87:chipyard.TestHarness.RocketConfig.fir@101436.4]
  assign _T_817 = setMatches[0] & abc_mshrs_0_io_status_bits_nestC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101099.4]
  assign _T_818 = setMatches[1] & abc_mshrs_1_io_status_bits_nestC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101100.4]
  assign _T_824 = _T_817 | _T_818; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101106.4]
  assign _T_819 = setMatches[2] & abc_mshrs_2_io_status_bits_nestC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101101.4]
  assign _T_825 = _T_824 | _T_819; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101107.4]
  assign _T_820 = setMatches[3] & abc_mshrs_3_io_status_bits_nestC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101102.4]
  assign _T_826 = _T_825 | _T_820; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101108.4]
  assign _T_821 = setMatches[4] & abc_mshrs_4_io_status_bits_nestC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101103.4]
  assign _T_827 = _T_826 | _T_821; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101109.4]
  assign _T_822 = setMatches[5] & bc_mshr_io_status_bits_nestC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101104.4]
  assign _T_828 = _T_827 | _T_822; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101110.4]
  assign _T_823 = setMatches[6] & c_mshr_io_status_bits_nestC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101105.4]
  assign _T_829 = _T_828 | _T_823; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101111.4]
  assign nestC = _T_829 & request_bits_prio_2; // @[Scheduler.scala 169:70:chipyard.TestHarness.RocketConfig.fir@101114.4]
  assign _T_1083 = nestC & _T_1072; // @[Scheduler.scala 249:13:chipyard.TestHarness.RocketConfig.fir@101440.4]
  assign _T_1085 = _T_1083 & _T_1079; // @[Scheduler.scala 249:56:chipyard.TestHarness.RocketConfig.fir@101442.4]
  assign request_alloc_cases = _T_1074 | _T_1085; // @[Scheduler.scala 248:112:chipyard.TestHarness.RocketConfig.fir@101443.4]
  assign lowerMatches = setMatches & prioFilter; // @[Scheduler.scala 172:33:chipyard.TestHarness.RocketConfig.fir@101119.4]
  assign _T_834 = |lowerMatches; // @[Scheduler.scala 174:31:chipyard.TestHarness.RocketConfig.fir@101120.4]
  assign _T_837 = ~nestC; // @[Scheduler.scala 174:47:chipyard.TestHarness.RocketConfig.fir@101123.4]
  assign _T_838 = _T_834 & _T_837; // @[Scheduler.scala 174:44:chipyard.TestHarness.RocketConfig.fir@101124.4]
  assign _T_775 = setMatches[0] & abc_mshrs_0_io_status_bits_blockC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101053.4]
  assign _T_776 = setMatches[1] & abc_mshrs_1_io_status_bits_blockC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101054.4]
  assign _T_782 = _T_775 | _T_776; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101060.4]
  assign _T_777 = setMatches[2] & abc_mshrs_2_io_status_bits_blockC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101055.4]
  assign _T_783 = _T_782 | _T_777; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101061.4]
  assign _T_778 = setMatches[3] & abc_mshrs_3_io_status_bits_blockC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101056.4]
  assign _T_784 = _T_783 | _T_778; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101062.4]
  assign _T_779 = setMatches[4] & abc_mshrs_4_io_status_bits_blockC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101057.4]
  assign _T_785 = _T_784 | _T_779; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101063.4]
  assign _T_780 = setMatches[5] & bc_mshr_io_status_bits_blockC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101058.4]
  assign _T_786 = _T_785 | _T_780; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101064.4]
  assign _T_781 = setMatches[6] & c_mshr_io_status_bits_blockC; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101059.4]
  assign _T_787 = _T_786 | _T_781; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101065.4]
  assign blockC = _T_787 & request_bits_prio_2; // @[Scheduler.scala 165:70:chipyard.TestHarness.RocketConfig.fir@101068.4]
  assign _T_841 = ~blockC; // @[Scheduler.scala 174:68:chipyard.TestHarness.RocketConfig.fir@101127.4]
  assign queue = _T_838 & _T_841; // @[Scheduler.scala 174:65:chipyard.TestHarness.RocketConfig.fir@101128.4]
  assign _T_847 = lowerMatches[5] ? 7'h20 : lowerMatches; // @[Scheduler.scala 190:8:chipyard.TestHarness.RocketConfig.fir@101134.4]
  assign lowerMatches1 = lowerMatches[6] ? 7'h40 : _T_847; // @[Scheduler.scala 189:8:chipyard.TestHarness.RocketConfig.fir@101135.4]
  assign _T_853 = mshr_selectOH & lowerMatches1; // @[Scheduler.scala 199:38:chipyard.TestHarness.RocketConfig.fir@101145.4]
  assign _T_854 = |_T_853; // @[Scheduler.scala 199:58:chipyard.TestHarness.RocketConfig.fir@101146.4]
  assign _T_855 = c_pop | request_bits_prio_2; // @[Scheduler.scala 200:33:chipyard.TestHarness.RocketConfig.fir@101147.4]
  assign _T_856 = ~c_pop; // @[Scheduler.scala 200:58:chipyard.TestHarness.RocketConfig.fir@101148.4]
  assign _T_858 = ~b_pop; // @[Scheduler.scala 200:101:chipyard.TestHarness.RocketConfig.fir@101150.4]
  assign _T_859 = ~a_pop; // @[Scheduler.scala 200:109:chipyard.TestHarness.RocketConfig.fir@101151.4]
  assign _T_860 = b_pop ? _T_858 : _T_859; // @[Scheduler.scala 200:69:chipyard.TestHarness.RocketConfig.fir@101152.4]
  assign _T_861 = _T_855 ? _T_856 : _T_860; // @[Scheduler.scala 200:26:chipyard.TestHarness.RocketConfig.fir@101153.4]
  assign bypassMatches = _T_854 & _T_861; // @[Scheduler.scala 199:61:chipyard.TestHarness.RocketConfig.fir@101154.4]
  assign bypassQueue = schedule_reload & bypassMatches; // @[Scheduler.scala 245:37:chipyard.TestHarness.RocketConfig.fir@101428.4]
  assign _T_1086 = bypassQueue | requests_io_push_ready; // @[Scheduler.scala 250:66:chipyard.TestHarness.RocketConfig.fir@101444.4]
  assign _T_1087 = queue & _T_1086; // @[Scheduler.scala 250:50:chipyard.TestHarness.RocketConfig.fir@101445.4]
  assign request_ready = request_alloc_cases | _T_1087; // @[Scheduler.scala 250:40:chipyard.TestHarness.RocketConfig.fir@101446.4]
  assign _T_718 = directory_io_ready & request_ready; // @[Scheduler.scala 156:44:chipyard.TestHarness.RocketConfig.fir@100989.4]
  assign _T_720 = ~sinkC_io_req_valid; // @[Scheduler.scala 157:64:chipyard.TestHarness.RocketConfig.fir@100992.4]
  assign _T_721 = _T_718 & _T_720; // @[Scheduler.scala 157:61:chipyard.TestHarness.RocketConfig.fir@100993.4]
  assign _T_725 = ~sinkX_io_req_valid; // @[Scheduler.scala 158:87:chipyard.TestHarness.RocketConfig.fir@100998.4]
  assign _T_843 = request_valid & nestC; // @[Scheduler.scala 182:33:chipyard.TestHarness.RocketConfig.fir@101130.4]
  assign _T_844 = request_valid & queue; // @[Scheduler.scala 184:31:chipyard.TestHarness.RocketConfig.fir@101131.4]
  assign bypass = _T_844 & bypassMatches; // @[Scheduler.scala 202:39:chipyard.TestHarness.RocketConfig.fir@101158.4]
  assign _T_864 = may_pop | bypass; // @[Scheduler.scala 203:49:chipyard.TestHarness.RocketConfig.fir@101159.4]
  assign will_reload = schedule_reload & _T_864; // @[Scheduler.scala 203:37:chipyard.TestHarness.RocketConfig.fir@101160.4]
  assign _T_866 = ~bypass; // @[Scheduler.scala 204:48:chipyard.TestHarness.RocketConfig.fir@101162.4]
  assign will_pop = _T_1062 & _T_866; // @[Scheduler.scala 204:45:chipyard.TestHarness.RocketConfig.fir@101163.4]
  assign _T_878 = requests_io_valid[14] | request_bits_prio_2; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101176.4]
  assign _T_879 = ~requests_io_valid[14]; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101177.4]
  assign _T_881 = ~requests_io_valid[7]; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101179.4]
  assign _T_882 = ~requests_io_valid[0]; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101180.4]
  assign _T_883 = requests_io_valid[7] ? _T_881 : _T_882; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101181.4]
  assign _T_884 = _T_878 ? _T_879 : _T_883; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101182.4]
  assign _T_885 = lowerMatches1[0] & _T_884; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101183.4]
  assign _T_886 = requests_io_valid[0] | requests_io_valid[7]; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101184.4]
  assign _T_887 = _T_886 | requests_io_valid[14]; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101185.4]
  assign _T_889 = _T_844 & _T_885; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101187.4]
  assign _T_890 = _T_887 | _T_889; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101188.4]
  assign _T_891 = abc_mshrs_0_io_schedule_bits_reload & _T_890; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101189.4]
  assign _T_893_prio_0 = _T_889 ? request_bits_prio_0 : requests_io_data_prio_0; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  assign _T_893_prio_1 = _T_889 ? 1'h0 : requests_io_data_prio_1; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  assign _T_893_prio_2 = _T_889 ? request_bits_prio_2 : requests_io_data_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  assign _T_893_control = _T_889 ? request_bits_control : requests_io_data_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  assign _T_893_opcode = _T_889 ? request_bits_opcode : requests_io_data_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  assign _T_893_param = _T_889 ? request_bits_param : requests_io_data_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  assign _T_893_size = _T_889 ? request_bits_size : requests_io_data_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  assign _T_893_source = _T_889 ? request_bits_source : requests_io_data_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  assign _T_893_tag = _T_889 ? request_bits_tag : requests_io_data_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  assign _T_893_offset = _T_889 ? request_bits_offset : requests_io_data_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  assign _T_893_put = _T_889 ? request_bits_put : requests_io_data_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101193.4]
  assign _T_894 = abc_mshrs_0_io_allocate_bits_tag == abc_mshrs_0_io_status_bits_tag; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101196.4]
  assign _T_895 = mshr_selectOH[0] & _T_891; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101198.4]
  assign _T_901 = requests_io_valid[15] | request_bits_prio_2; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101206.4]
  assign _T_902 = ~requests_io_valid[15]; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101207.4]
  assign _T_904 = ~requests_io_valid[8]; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101209.4]
  assign _T_905 = ~requests_io_valid[1]; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101210.4]
  assign _T_906 = requests_io_valid[8] ? _T_904 : _T_905; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101211.4]
  assign _T_907 = _T_901 ? _T_902 : _T_906; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101212.4]
  assign _T_908 = lowerMatches1[1] & _T_907; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101213.4]
  assign _T_909 = requests_io_valid[1] | requests_io_valid[8]; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101214.4]
  assign _T_910 = _T_909 | requests_io_valid[15]; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101215.4]
  assign _T_912 = _T_844 & _T_908; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101217.4]
  assign _T_913 = _T_910 | _T_912; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101218.4]
  assign _T_914 = abc_mshrs_1_io_schedule_bits_reload & _T_913; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101219.4]
  assign _T_916_prio_0 = _T_912 ? request_bits_prio_0 : requests_io_data_prio_0; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  assign _T_916_prio_1 = _T_912 ? 1'h0 : requests_io_data_prio_1; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  assign _T_916_prio_2 = _T_912 ? request_bits_prio_2 : requests_io_data_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  assign _T_916_control = _T_912 ? request_bits_control : requests_io_data_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  assign _T_916_opcode = _T_912 ? request_bits_opcode : requests_io_data_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  assign _T_916_param = _T_912 ? request_bits_param : requests_io_data_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  assign _T_916_size = _T_912 ? request_bits_size : requests_io_data_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  assign _T_916_source = _T_912 ? request_bits_source : requests_io_data_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  assign _T_916_tag = _T_912 ? request_bits_tag : requests_io_data_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  assign _T_916_offset = _T_912 ? request_bits_offset : requests_io_data_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  assign _T_916_put = _T_912 ? request_bits_put : requests_io_data_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101223.4]
  assign _T_917 = abc_mshrs_1_io_allocate_bits_tag == abc_mshrs_1_io_status_bits_tag; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101226.4]
  assign _T_918 = mshr_selectOH[1] & _T_914; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101228.4]
  assign _T_924 = requests_io_valid[16] | request_bits_prio_2; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101236.4]
  assign _T_925 = ~requests_io_valid[16]; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101237.4]
  assign _T_927 = ~requests_io_valid[9]; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101239.4]
  assign _T_928 = ~requests_io_valid[2]; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101240.4]
  assign _T_929 = requests_io_valid[9] ? _T_927 : _T_928; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101241.4]
  assign _T_930 = _T_924 ? _T_925 : _T_929; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101242.4]
  assign _T_931 = lowerMatches1[2] & _T_930; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101243.4]
  assign _T_932 = requests_io_valid[2] | requests_io_valid[9]; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101244.4]
  assign _T_933 = _T_932 | requests_io_valid[16]; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101245.4]
  assign _T_935 = _T_844 & _T_931; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101247.4]
  assign _T_936 = _T_933 | _T_935; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101248.4]
  assign _T_937 = abc_mshrs_2_io_schedule_bits_reload & _T_936; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101249.4]
  assign _T_939_prio_0 = _T_935 ? request_bits_prio_0 : requests_io_data_prio_0; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  assign _T_939_prio_1 = _T_935 ? 1'h0 : requests_io_data_prio_1; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  assign _T_939_prio_2 = _T_935 ? request_bits_prio_2 : requests_io_data_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  assign _T_939_control = _T_935 ? request_bits_control : requests_io_data_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  assign _T_939_opcode = _T_935 ? request_bits_opcode : requests_io_data_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  assign _T_939_param = _T_935 ? request_bits_param : requests_io_data_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  assign _T_939_size = _T_935 ? request_bits_size : requests_io_data_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  assign _T_939_source = _T_935 ? request_bits_source : requests_io_data_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  assign _T_939_tag = _T_935 ? request_bits_tag : requests_io_data_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  assign _T_939_offset = _T_935 ? request_bits_offset : requests_io_data_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  assign _T_939_put = _T_935 ? request_bits_put : requests_io_data_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101253.4]
  assign _T_940 = abc_mshrs_2_io_allocate_bits_tag == abc_mshrs_2_io_status_bits_tag; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101256.4]
  assign _T_941 = mshr_selectOH[2] & _T_937; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101258.4]
  assign _T_947 = requests_io_valid[17] | request_bits_prio_2; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101266.4]
  assign _T_948 = ~requests_io_valid[17]; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101267.4]
  assign _T_950 = ~requests_io_valid[10]; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101269.4]
  assign _T_951 = ~requests_io_valid[3]; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101270.4]
  assign _T_952 = requests_io_valid[10] ? _T_950 : _T_951; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101271.4]
  assign _T_953 = _T_947 ? _T_948 : _T_952; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101272.4]
  assign _T_954 = lowerMatches1[3] & _T_953; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101273.4]
  assign _T_955 = requests_io_valid[3] | requests_io_valid[10]; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101274.4]
  assign _T_956 = _T_955 | requests_io_valid[17]; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101275.4]
  assign _T_958 = _T_844 & _T_954; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101277.4]
  assign _T_959 = _T_956 | _T_958; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101278.4]
  assign _T_960 = abc_mshrs_3_io_schedule_bits_reload & _T_959; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101279.4]
  assign _T_962_prio_0 = _T_958 ? request_bits_prio_0 : requests_io_data_prio_0; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  assign _T_962_prio_1 = _T_958 ? 1'h0 : requests_io_data_prio_1; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  assign _T_962_prio_2 = _T_958 ? request_bits_prio_2 : requests_io_data_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  assign _T_962_control = _T_958 ? request_bits_control : requests_io_data_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  assign _T_962_opcode = _T_958 ? request_bits_opcode : requests_io_data_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  assign _T_962_param = _T_958 ? request_bits_param : requests_io_data_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  assign _T_962_size = _T_958 ? request_bits_size : requests_io_data_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  assign _T_962_source = _T_958 ? request_bits_source : requests_io_data_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  assign _T_962_tag = _T_958 ? request_bits_tag : requests_io_data_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  assign _T_962_offset = _T_958 ? request_bits_offset : requests_io_data_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  assign _T_962_put = _T_958 ? request_bits_put : requests_io_data_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101283.4]
  assign _T_963 = abc_mshrs_3_io_allocate_bits_tag == abc_mshrs_3_io_status_bits_tag; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101286.4]
  assign _T_964 = mshr_selectOH[3] & _T_960; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101288.4]
  assign _T_970 = requests_io_valid[18] | request_bits_prio_2; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101296.4]
  assign _T_971 = ~requests_io_valid[18]; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101297.4]
  assign _T_973 = ~requests_io_valid[11]; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101299.4]
  assign _T_974 = ~requests_io_valid[4]; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101300.4]
  assign _T_975 = requests_io_valid[11] ? _T_973 : _T_974; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101301.4]
  assign _T_976 = _T_970 ? _T_971 : _T_975; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101302.4]
  assign _T_977 = lowerMatches1[4] & _T_976; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101303.4]
  assign _T_978 = requests_io_valid[4] | requests_io_valid[11]; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101304.4]
  assign _T_979 = _T_978 | requests_io_valid[18]; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101305.4]
  assign _T_981 = _T_844 & _T_977; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101307.4]
  assign _T_982 = _T_979 | _T_981; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101308.4]
  assign _T_983 = abc_mshrs_4_io_schedule_bits_reload & _T_982; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101309.4]
  assign _T_985_prio_0 = _T_981 ? request_bits_prio_0 : requests_io_data_prio_0; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  assign _T_985_prio_1 = _T_981 ? 1'h0 : requests_io_data_prio_1; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  assign _T_985_prio_2 = _T_981 ? request_bits_prio_2 : requests_io_data_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  assign _T_985_control = _T_981 ? request_bits_control : requests_io_data_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  assign _T_985_opcode = _T_981 ? request_bits_opcode : requests_io_data_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  assign _T_985_param = _T_981 ? request_bits_param : requests_io_data_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  assign _T_985_size = _T_981 ? request_bits_size : requests_io_data_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  assign _T_985_source = _T_981 ? request_bits_source : requests_io_data_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  assign _T_985_tag = _T_981 ? request_bits_tag : requests_io_data_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  assign _T_985_offset = _T_981 ? request_bits_offset : requests_io_data_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  assign _T_985_put = _T_981 ? request_bits_put : requests_io_data_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101313.4]
  assign _T_986 = abc_mshrs_4_io_allocate_bits_tag == abc_mshrs_4_io_status_bits_tag; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101316.4]
  assign _T_987 = mshr_selectOH[4] & _T_983; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101318.4]
  assign _T_993 = requests_io_valid[19] | request_bits_prio_2; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101326.4]
  assign _T_994 = ~requests_io_valid[19]; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101327.4]
  assign _T_996 = ~requests_io_valid[12]; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101329.4]
  assign _T_997 = ~requests_io_valid[5]; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101330.4]
  assign _T_998 = requests_io_valid[12] ? _T_996 : _T_997; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101331.4]
  assign _T_999 = _T_993 ? _T_994 : _T_998; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101332.4]
  assign _T_1000 = lowerMatches1[5] & _T_999; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101333.4]
  assign _T_1001 = requests_io_valid[5] | requests_io_valid[12]; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101334.4]
  assign _T_1002 = _T_1001 | requests_io_valid[19]; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101335.4]
  assign _T_1004 = _T_844 & _T_1000; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101337.4]
  assign _T_1005 = _T_1002 | _T_1004; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101338.4]
  assign _T_1006 = bc_mshr_io_schedule_bits_reload & _T_1005; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101339.4]
  assign _T_1008_prio_1 = _T_1004 ? 1'h0 : requests_io_data_prio_1; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  assign _T_1008_prio_2 = _T_1004 ? request_bits_prio_2 : requests_io_data_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  assign _T_1008_control = _T_1004 ? request_bits_control : requests_io_data_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  assign _T_1008_opcode = _T_1004 ? request_bits_opcode : requests_io_data_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  assign _T_1008_param = _T_1004 ? request_bits_param : requests_io_data_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  assign _T_1008_size = _T_1004 ? request_bits_size : requests_io_data_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  assign _T_1008_source = _T_1004 ? request_bits_source : requests_io_data_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  assign _T_1008_tag = _T_1004 ? request_bits_tag : requests_io_data_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  assign _T_1008_offset = _T_1004 ? request_bits_offset : requests_io_data_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  assign _T_1008_put = _T_1004 ? request_bits_put : requests_io_data_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101343.4]
  assign _T_1009 = bc_mshr_io_allocate_bits_tag == bc_mshr_io_status_bits_tag; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101346.4]
  assign _T_1010 = mshr_selectOH[5] & _T_1006; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101348.4]
  assign _T_1016 = requests_io_valid[20] | request_bits_prio_2; // @[Scheduler.scala 218:35:chipyard.TestHarness.RocketConfig.fir@101356.4]
  assign _T_1017 = ~requests_io_valid[20]; // @[Scheduler.scala 218:60:chipyard.TestHarness.RocketConfig.fir@101357.4]
  assign _T_1019 = ~requests_io_valid[13]; // @[Scheduler.scala 218:103:chipyard.TestHarness.RocketConfig.fir@101359.4]
  assign _T_1020 = ~requests_io_valid[6]; // @[Scheduler.scala 218:111:chipyard.TestHarness.RocketConfig.fir@101360.4]
  assign _T_1021 = requests_io_valid[13] ? _T_1019 : _T_1020; // @[Scheduler.scala 218:71:chipyard.TestHarness.RocketConfig.fir@101361.4]
  assign _T_1022 = _T_1016 ? _T_1017 : _T_1021; // @[Scheduler.scala 218:28:chipyard.TestHarness.RocketConfig.fir@101362.4]
  assign _T_1023 = lowerMatches1[6] & _T_1022; // @[Scheduler.scala 217:42:chipyard.TestHarness.RocketConfig.fir@101363.4]
  assign _T_1024 = requests_io_valid[6] | requests_io_valid[13]; // @[Scheduler.scala 219:25:chipyard.TestHarness.RocketConfig.fir@101364.4]
  assign _T_1025 = _T_1024 | requests_io_valid[20]; // @[Scheduler.scala 219:34:chipyard.TestHarness.RocketConfig.fir@101365.4]
  assign _T_1027 = _T_844 & _T_1023; // @[Scheduler.scala 220:41:chipyard.TestHarness.RocketConfig.fir@101367.4]
  assign _T_1028 = _T_1025 | _T_1027; // @[Scheduler.scala 221:61:chipyard.TestHarness.RocketConfig.fir@101368.4]
  assign _T_1029 = c_mshr_io_schedule_bits_reload & _T_1028; // @[Scheduler.scala 221:49:chipyard.TestHarness.RocketConfig.fir@101369.4]
  assign _T_1031_prio_2 = _T_1027 ? request_bits_prio_2 : requests_io_data_prio_2; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  assign _T_1031_control = _T_1027 ? request_bits_control : requests_io_data_control; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  assign _T_1031_opcode = _T_1027 ? request_bits_opcode : requests_io_data_opcode; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  assign _T_1031_param = _T_1027 ? request_bits_param : requests_io_data_param; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  assign _T_1031_size = _T_1027 ? request_bits_size : requests_io_data_size; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  assign _T_1031_source = _T_1027 ? request_bits_source : requests_io_data_source; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  assign _T_1031_tag = _T_1027 ? request_bits_tag : requests_io_data_tag; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  assign _T_1031_offset = _T_1027 ? request_bits_offset : requests_io_data_offset; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  assign _T_1031_put = _T_1027 ? request_bits_put : requests_io_data_put; // @[Scheduler.scala 222:30:chipyard.TestHarness.RocketConfig.fir@101373.4]
  assign _T_1032 = c_mshr_io_allocate_bits_tag == c_mshr_io_status_bits_tag; // @[Scheduler.scala 224:57:chipyard.TestHarness.RocketConfig.fir@101376.4]
  assign _T_1033 = mshr_selectOH[6] & _T_1029; // @[Scheduler.scala 225:32:chipyard.TestHarness.RocketConfig.fir@101378.4]
  assign _T_1034 = ~requests_io_valid; // @[Scheduler.scala 229:25:chipyard.TestHarness.RocketConfig.fir@101380.4]
  assign _GEN_146 = {{7'd0}, requests_io_valid[20:7]}; // @[Scheduler.scala 229:44:chipyard.TestHarness.RocketConfig.fir@101382.4]
  assign _T_1036 = _T_1034 | _GEN_146; // @[Scheduler.scala 229:44:chipyard.TestHarness.RocketConfig.fir@101382.4]
  assign _GEN_147 = {{14'd0}, requests_io_valid[20:14]}; // @[Scheduler.scala 229:82:chipyard.TestHarness.RocketConfig.fir@101384.4]
  assign _T_1038 = _T_1036 | _GEN_147; // @[Scheduler.scala 229:82:chipyard.TestHarness.RocketConfig.fir@101384.4]
  assign prio_requests = ~_T_1038; // @[Scheduler.scala 229:23:chipyard.TestHarness.RocketConfig.fir@101385.4]
  assign _T_1041 = _T_849 & prio_requests; // @[Scheduler.scala 230:77:chipyard.TestHarness.RocketConfig.fir@101388.4]
  assign _T_1044 = |_T_1041[20:16]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101391.4]
  assign _GEN_148 = {{11'd0}, _T_1041[20:16]}; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101392.4]
  assign _T_1045 = _GEN_148 | _T_1041[15:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101392.4]
  assign _T_1048 = |_T_1045[15:8]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101395.4]
  assign _T_1049 = _T_1045[15:8] | _T_1045[7:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101396.4]
  assign _T_1052 = |_T_1049[7:4]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101399.4]
  assign _T_1053 = _T_1049[7:4] | _T_1049[3:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101400.4]
  assign _T_1056 = |_T_1053[3:2]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101403.4]
  assign _T_1057 = _T_1053[3:2] | _T_1053[1:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101404.4]
  assign _T_1061 = {_T_1048,_T_1052,_T_1056,_T_1057[1]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101408.4]
  assign mshr_uses_directory_for_lb = will_pop & lb_tag_mismatch; // @[Scheduler.scala 237:45:chipyard.TestHarness.RocketConfig.fir@101415.4]
  assign _T_1063 = bypass ? request_bits_tag : requests_io_data_tag; // @[Scheduler.scala 238:63:chipyard.TestHarness.RocketConfig.fir@101416.4]
  assign _T_1064 = scheduleTag != _T_1063; // @[Scheduler.scala 238:56:chipyard.TestHarness.RocketConfig.fir@101417.4]
  assign mshr_uses_directory = will_reload & _T_1064; // @[Scheduler.scala 238:41:chipyard.TestHarness.RocketConfig.fir@101418.4]
  assign alloc_uses_directory = request_valid & request_alloc_cases; // @[Scheduler.scala 251:44:chipyard.TestHarness.RocketConfig.fir@101448.4]
  assign _T_1093 = ~bypassQueue; // @[Scheduler.scala 259:55:chipyard.TestHarness.RocketConfig.fir@101456.4]
  assign _T_1098 = |lowerMatches1[6:4]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101463.4]
  assign _GEN_149 = {{1'd0}, lowerMatches1[6:4]}; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101464.4]
  assign _T_1099 = _GEN_149 | lowerMatches1[3:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101464.4]
  assign _T_1102 = |_T_1099[3:2]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101467.4]
  assign _T_1103 = _T_1099[3:2] | _T_1099[1:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101468.4]
  assign _T_1106 = {_T_1098,_T_1102,_T_1103[1]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101471.4]
  assign _T_1124 = {lowerMatches1, 14'h0}; // @[Scheduler.scala 265:30:chipyard.TestHarness.RocketConfig.fir@101489.4]
  assign _T_1127 = |_T_1124[20:16]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101492.4]
  assign _GEN_151 = {{11'd0}, _T_1124[20:16]}; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101493.4]
  assign _T_1128 = _GEN_151 | _T_1124[15:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101493.4]
  assign _T_1131 = |_T_1128[15:8]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101496.4]
  assign _T_1132 = _T_1128[15:8] | _T_1128[7:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101497.4]
  assign _T_1135 = |_T_1132[7:4]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101500.4]
  assign _T_1136 = _T_1132[7:4] | _T_1132[3:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101501.4]
  assign _T_1139 = |_T_1136[3:2]; // @[OneHot.scala 32:14:chipyard.TestHarness.RocketConfig.fir@101504.4]
  assign _T_1140 = _T_1136[3:2] | _T_1136[1:0]; // @[OneHot.scala 32:28:chipyard.TestHarness.RocketConfig.fir@101505.4]
  assign _T_1145 = {_T_1127,_T_1131,_T_1135,_T_1139,_T_1140[1]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@101510.4]
  assign _T_1146 = request_bits_prio_0 ? _T_1106 : 3'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101511.4]
  assign _T_1148 = request_bits_prio_2 ? _T_1145 : 5'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101513.4]
  assign _T_1149 = {{1'd0}, _T_1146}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101514.4]
  assign _GEN_152 = {{1'd0}, _T_1149}; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101515.4]
  assign _T_1153 = {_T_1070, 1'h0}; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@101520.4]
  assign _T_1155 = _T_1070 | _T_1153[6:0]; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@101522.4]
  assign _T_1156 = {_T_1155, 2'h0}; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@101523.4]
  assign _T_1158 = _T_1155 | _T_1156[6:0]; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@101525.4]
  assign _T_1159 = {_T_1158, 4'h0}; // @[package.scala 199:48:chipyard.TestHarness.RocketConfig.fir@101526.4]
  assign _T_1161 = _T_1158 | _T_1159[6:0]; // @[package.scala 199:43:chipyard.TestHarness.RocketConfig.fir@101528.4]
  assign _T_1163 = {_T_1161, 1'h0}; // @[Scheduler.scala 267:47:chipyard.TestHarness.RocketConfig.fir@101530.4]
  assign _T_1164 = ~_T_1163; // @[Scheduler.scala 267:23:chipyard.TestHarness.RocketConfig.fir@101531.4]
  assign _GEN_153 = {{1'd0}, _T_1070}; // @[Scheduler.scala 267:53:chipyard.TestHarness.RocketConfig.fir@101533.4]
  assign _T_1166 = _T_1164 & _GEN_153; // @[Scheduler.scala 267:53:chipyard.TestHarness.RocketConfig.fir@101533.4]
  assign _GEN_154 = {{1'd0}, prioFilter}; // @[Scheduler.scala 267:69:chipyard.TestHarness.RocketConfig.fir@101534.4]
  assign mshr_insertOH = _T_1166 & _GEN_154; // @[Scheduler.scala 267:69:chipyard.TestHarness.RocketConfig.fir@101534.4]
  assign _T_1175 = request_valid & alloc; // @[Scheduler.scala 269:25:chipyard.TestHarness.RocketConfig.fir@101543.4]
  assign _T_1176 = _T_1175 & mshr_insertOH[0]; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101544.4]
  assign _T_1178 = _T_1176 & _T_1072; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101546.4]
  assign _T_1180 = _T_1175 & mshr_insertOH[1]; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101553.4]
  assign _T_1182 = _T_1180 & _T_1072; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101555.4]
  assign _T_1184 = _T_1175 & mshr_insertOH[2]; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101562.4]
  assign _T_1186 = _T_1184 & _T_1072; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101564.4]
  assign _T_1188 = _T_1175 & mshr_insertOH[3]; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101571.4]
  assign _T_1190 = _T_1188 & _T_1072; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101573.4]
  assign _T_1192 = _T_1175 & mshr_insertOH[4]; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101580.4]
  assign _T_1194 = _T_1192 & _T_1072; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101582.4]
  assign _T_1196 = _T_1175 & mshr_insertOH[5]; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101589.4]
  assign _T_1198 = _T_1196 & _T_1072; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101591.4]
  assign _T_1200 = _T_1175 & mshr_insertOH[6]; // @[Scheduler.scala 269:34:chipyard.TestHarness.RocketConfig.fir@101598.4]
  assign _T_1202 = _T_1200 & _T_1072; // @[Scheduler.scala 269:39:chipyard.TestHarness.RocketConfig.fir@101600.4]
  assign _GEN_85 = _T_1202 | _T_1033; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  assign _GEN_88 = _T_1202 ? request_bits_prio_2 : _T_1031_prio_2; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  assign _GEN_89 = _T_1202 ? request_bits_control : _T_1031_control; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  assign _GEN_90 = _T_1202 ? request_bits_opcode : _T_1031_opcode; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  assign _GEN_91 = _T_1202 ? request_bits_param : _T_1031_param; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  assign _GEN_92 = _T_1202 ? request_bits_size : _T_1031_size; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  assign _GEN_93 = _T_1202 ? request_bits_source : _T_1031_source; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  assign _GEN_94 = _T_1202 ? request_bits_tag : _T_1031_tag; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  assign _GEN_95 = _T_1202 ? request_bits_offset : _T_1031_offset; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  assign _GEN_96 = _T_1202 ? request_bits_put : _T_1031_put; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  assign _GEN_97 = _T_1202 ? request_bits_set : c_mshr_io_status_bits_set; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  assign _GEN_98 = _T_1202 ? 1'h0 : _T_1032; // @[Scheduler.scala 269:83:chipyard.TestHarness.RocketConfig.fir@101601.4]
  assign _T_1212 = _T_831 | reset; // @[Scheduler.scala 280:12:chipyard.TestHarness.RocketConfig.fir@101619.6]
  assign _T_1213 = ~_T_1212; // @[Scheduler.scala 280:12:chipyard.TestHarness.RocketConfig.fir@101620.6]
  assign _T_1216 = _T_843 & _T_1079; // @[Scheduler.scala 284:32:chipyard.TestHarness.RocketConfig.fir@101629.4]
  assign _T_1218 = _T_1216 & _T_1072; // @[Scheduler.scala 284:59:chipyard.TestHarness.RocketConfig.fir@101631.4]
  assign _T_1237 = bc_mshr_io_status_bits_set == sinkC_io_set; // @[Scheduler.scala 304:63:chipyard.TestHarness.RocketConfig.fir@101682.4]
  assign _T_1238 = bc_mshr_io_status_valid & _T_1237; // @[Scheduler.scala 304:33:chipyard.TestHarness.RocketConfig.fir@101683.4]
  assign _T_1239 = abc_mshrs_0_io_status_bits_set == sinkC_io_set; // @[Scheduler.scala 306:74:chipyard.TestHarness.RocketConfig.fir@101684.4]
  assign _T_1240 = abc_mshrs_0_io_status_valid & _T_1239; // @[Scheduler.scala 306:50:chipyard.TestHarness.RocketConfig.fir@101685.4]
  assign _T_1241 = abc_mshrs_1_io_status_bits_set == sinkC_io_set; // @[Scheduler.scala 306:74:chipyard.TestHarness.RocketConfig.fir@101686.4]
  assign _T_1242 = abc_mshrs_1_io_status_valid & _T_1241; // @[Scheduler.scala 306:50:chipyard.TestHarness.RocketConfig.fir@101687.4]
  assign _T_1243 = abc_mshrs_2_io_status_bits_set == sinkC_io_set; // @[Scheduler.scala 306:74:chipyard.TestHarness.RocketConfig.fir@101688.4]
  assign _T_1244 = abc_mshrs_2_io_status_valid & _T_1243; // @[Scheduler.scala 306:50:chipyard.TestHarness.RocketConfig.fir@101689.4]
  assign _T_1245 = abc_mshrs_3_io_status_bits_set == sinkC_io_set; // @[Scheduler.scala 306:74:chipyard.TestHarness.RocketConfig.fir@101690.4]
  assign _T_1246 = abc_mshrs_3_io_status_valid & _T_1245; // @[Scheduler.scala 306:50:chipyard.TestHarness.RocketConfig.fir@101691.4]
  assign _T_1247 = abc_mshrs_4_io_status_bits_set == sinkC_io_set; // @[Scheduler.scala 306:74:chipyard.TestHarness.RocketConfig.fir@101692.4]
  assign _T_1248 = abc_mshrs_4_io_status_valid & _T_1247; // @[Scheduler.scala 306:50:chipyard.TestHarness.RocketConfig.fir@101693.4]
  assign _T_1249 = _T_1240 ? abc_mshrs_0_io_status_bits_way : 3'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101694.4]
  assign _T_1250 = _T_1242 ? abc_mshrs_1_io_status_bits_way : 3'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101695.4]
  assign _T_1251 = _T_1244 ? abc_mshrs_2_io_status_bits_way : 3'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101696.4]
  assign _T_1252 = _T_1246 ? abc_mshrs_3_io_status_bits_way : 3'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101697.4]
  assign _T_1253 = _T_1248 ? abc_mshrs_4_io_status_bits_way : 3'h0; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101698.4]
  assign _T_1254 = _T_1249 | _T_1250; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101699.4]
  assign _T_1255 = _T_1254 | _T_1251; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101700.4]
  assign _T_1256 = _T_1255 | _T_1252; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101701.4]
  assign _T_1257 = _T_1256 | _T_1253; // @[Mux.scala 27:72:chipyard.TestHarness.RocketConfig.fir@101702.4]
  assign _T_1260_0 = abc_mshrs_0_io_status_bits_way; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101709.4]
  assign _T_1260_1 = abc_mshrs_1_io_status_bits_way; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101710.4]
  assign _GEN_128 = 3'h1 == sinkD_io_source ? _T_1260_1 : _T_1260_0; // @[Scheduler.scala 308:16:chipyard.TestHarness.RocketConfig.fir@101716.4]
  assign _T_1260_2 = abc_mshrs_2_io_status_bits_way; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101711.4]
  assign _GEN_129 = 3'h2 == sinkD_io_source ? _T_1260_2 : _GEN_128; // @[Scheduler.scala 308:16:chipyard.TestHarness.RocketConfig.fir@101716.4]
  assign _T_1260_3 = abc_mshrs_3_io_status_bits_way; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101712.4]
  assign _GEN_130 = 3'h3 == sinkD_io_source ? _T_1260_3 : _GEN_129; // @[Scheduler.scala 308:16:chipyard.TestHarness.RocketConfig.fir@101716.4]
  assign _T_1260_4 = abc_mshrs_4_io_status_bits_way; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101713.4]
  assign _GEN_131 = 3'h4 == sinkD_io_source ? _T_1260_4 : _GEN_130; // @[Scheduler.scala 308:16:chipyard.TestHarness.RocketConfig.fir@101716.4]
  assign _T_1260_5 = bc_mshr_io_status_bits_way; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101714.4]
  assign _GEN_132 = 3'h5 == sinkD_io_source ? _T_1260_5 : _GEN_131; // @[Scheduler.scala 308:16:chipyard.TestHarness.RocketConfig.fir@101716.4]
  assign _T_1260_6 = c_mshr_io_status_bits_way; // @[Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101707.4 Scheduler.scala 308:22:chipyard.TestHarness.RocketConfig.fir@101715.4]
  assign _T_1261_0 = abc_mshrs_0_io_status_bits_set; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101719.4]
  assign _T_1261_1 = abc_mshrs_1_io_status_bits_set; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101720.4]
  assign _GEN_135 = 3'h1 == sinkD_io_source ? _T_1261_1 : _T_1261_0; // @[Scheduler.scala 309:16:chipyard.TestHarness.RocketConfig.fir@101726.4]
  assign _T_1261_2 = abc_mshrs_2_io_status_bits_set; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101721.4]
  assign _GEN_136 = 3'h2 == sinkD_io_source ? _T_1261_2 : _GEN_135; // @[Scheduler.scala 309:16:chipyard.TestHarness.RocketConfig.fir@101726.4]
  assign _T_1261_3 = abc_mshrs_3_io_status_bits_set; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101722.4]
  assign _GEN_137 = 3'h3 == sinkD_io_source ? _T_1261_3 : _GEN_136; // @[Scheduler.scala 309:16:chipyard.TestHarness.RocketConfig.fir@101726.4]
  assign _T_1261_4 = abc_mshrs_4_io_status_bits_set; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101723.4]
  assign _GEN_138 = 3'h4 == sinkD_io_source ? _T_1261_4 : _GEN_137; // @[Scheduler.scala 309:16:chipyard.TestHarness.RocketConfig.fir@101726.4]
  assign _T_1261_5 = bc_mshr_io_status_bits_set; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101724.4]
  assign _GEN_139 = 3'h5 == sinkD_io_source ? _T_1261_5 : _GEN_138; // @[Scheduler.scala 309:16:chipyard.TestHarness.RocketConfig.fir@101726.4]
  assign _T_1261_6 = c_mshr_io_status_bits_set; // @[Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101717.4 Scheduler.scala 309:22:chipyard.TestHarness.RocketConfig.fir@101725.4]
  assign io_in_a_ready = sinkA_io_a_ready; // @[Scheduler.scala 58:14:chipyard.TestHarness.RocketConfig.fir@100079.4]
  assign io_in_b_valid = sourceB_io_b_valid; // @[Scheduler.scala 48:11:chipyard.TestHarness.RocketConfig.fir@100056.4]
  assign io_in_b_bits_param = sourceB_io_b_bits_param; // @[Scheduler.scala 48:11:chipyard.TestHarness.RocketConfig.fir@100056.4]
  assign io_in_b_bits_address = sourceB_io_b_bits_address; // @[Scheduler.scala 48:11:chipyard.TestHarness.RocketConfig.fir@100056.4]
  assign io_in_c_ready = sinkC_io_c_ready; // @[Scheduler.scala 59:14:chipyard.TestHarness.RocketConfig.fir@100080.4]
  assign io_in_d_valid = sourceD_io_d_valid; // @[Scheduler.scala 49:11:chipyard.TestHarness.RocketConfig.fir@100057.4]
  assign io_in_d_bits_opcode = sourceD_io_d_bits_opcode; // @[Scheduler.scala 49:11:chipyard.TestHarness.RocketConfig.fir@100057.4]
  assign io_in_d_bits_param = sourceD_io_d_bits_param; // @[Scheduler.scala 49:11:chipyard.TestHarness.RocketConfig.fir@100057.4]
  assign io_in_d_bits_size = sourceD_io_d_bits_size; // @[Scheduler.scala 49:11:chipyard.TestHarness.RocketConfig.fir@100057.4]
  assign io_in_d_bits_source = sourceD_io_d_bits_source; // @[Scheduler.scala 49:11:chipyard.TestHarness.RocketConfig.fir@100057.4]
  assign io_in_d_bits_sink = sourceD_io_d_bits_sink; // @[Scheduler.scala 49:11:chipyard.TestHarness.RocketConfig.fir@100057.4]
  assign io_in_d_bits_denied = sourceD_io_d_bits_denied; // @[Scheduler.scala 49:11:chipyard.TestHarness.RocketConfig.fir@100057.4]
  assign io_in_d_bits_data = sourceD_io_d_bits_data; // @[Scheduler.scala 49:11:chipyard.TestHarness.RocketConfig.fir@100057.4]
  assign io_in_d_bits_corrupt = sourceD_io_d_bits_corrupt; // @[Scheduler.scala 49:11:chipyard.TestHarness.RocketConfig.fir@100057.4]
  assign io_out_a_valid = sourceA_io_a_valid; // @[Scheduler.scala 45:12:chipyard.TestHarness.RocketConfig.fir@100053.4]
  assign io_out_a_bits_opcode = sourceA_io_a_bits_opcode; // @[Scheduler.scala 45:12:chipyard.TestHarness.RocketConfig.fir@100053.4]
  assign io_out_a_bits_param = sourceA_io_a_bits_param; // @[Scheduler.scala 45:12:chipyard.TestHarness.RocketConfig.fir@100053.4]
  assign io_out_a_bits_size = sourceA_io_a_bits_size; // @[Scheduler.scala 45:12:chipyard.TestHarness.RocketConfig.fir@100053.4]
  assign io_out_a_bits_source = sourceA_io_a_bits_source; // @[Scheduler.scala 45:12:chipyard.TestHarness.RocketConfig.fir@100053.4]
  assign io_out_a_bits_address = sourceA_io_a_bits_address; // @[Scheduler.scala 45:12:chipyard.TestHarness.RocketConfig.fir@100053.4]
  assign io_out_a_bits_mask = sourceA_io_a_bits_mask; // @[Scheduler.scala 45:12:chipyard.TestHarness.RocketConfig.fir@100053.4]
  assign io_out_a_bits_data = sourceA_io_a_bits_data; // @[Scheduler.scala 45:12:chipyard.TestHarness.RocketConfig.fir@100053.4]
  assign io_out_a_bits_corrupt = sourceA_io_a_bits_corrupt; // @[Scheduler.scala 45:12:chipyard.TestHarness.RocketConfig.fir@100053.4]
  assign io_out_c_valid = sourceC_io_c_valid; // @[Scheduler.scala 46:12:chipyard.TestHarness.RocketConfig.fir@100054.4]
  assign io_out_c_bits_opcode = sourceC_io_c_bits_opcode; // @[Scheduler.scala 46:12:chipyard.TestHarness.RocketConfig.fir@100054.4]
  assign io_out_c_bits_param = sourceC_io_c_bits_param; // @[Scheduler.scala 46:12:chipyard.TestHarness.RocketConfig.fir@100054.4]
  assign io_out_c_bits_size = sourceC_io_c_bits_size; // @[Scheduler.scala 46:12:chipyard.TestHarness.RocketConfig.fir@100054.4]
  assign io_out_c_bits_source = sourceC_io_c_bits_source; // @[Scheduler.scala 46:12:chipyard.TestHarness.RocketConfig.fir@100054.4]
  assign io_out_c_bits_address = sourceC_io_c_bits_address; // @[Scheduler.scala 46:12:chipyard.TestHarness.RocketConfig.fir@100054.4]
  assign io_out_c_bits_data = sourceC_io_c_bits_data; // @[Scheduler.scala 46:12:chipyard.TestHarness.RocketConfig.fir@100054.4]
  assign io_out_c_bits_corrupt = sourceC_io_c_bits_corrupt; // @[Scheduler.scala 46:12:chipyard.TestHarness.RocketConfig.fir@100054.4]
  assign io_out_d_ready = sinkD_io_d_ready; // @[Scheduler.scala 61:14:chipyard.TestHarness.RocketConfig.fir@100082.4]
  assign io_out_e_valid = sourceE_io_e_valid; // @[Scheduler.scala 47:12:chipyard.TestHarness.RocketConfig.fir@100055.4]
  assign io_out_e_bits_sink = sourceE_io_e_bits_sink; // @[Scheduler.scala 47:12:chipyard.TestHarness.RocketConfig.fir@100055.4]
  assign io_req_ready = sinkX_io_x_ready; // @[Scheduler.scala 62:14:chipyard.TestHarness.RocketConfig.fir@100083.4]
  assign io_resp_valid = sourceX_io_x_valid; // @[Scheduler.scala 50:11:chipyard.TestHarness.RocketConfig.fir@100058.4]
  assign sourceA_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100031.4]
  assign sourceA_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100032.4]
  assign sourceA_io_req_valid = _T_602[187]; // @[Scheduler.scala 133:18:chipyard.TestHarness.RocketConfig.fir@100954.4]
  assign sourceA_io_req_bits_tag = _T_602[186:175]; // @[Scheduler.scala 133:18:chipyard.TestHarness.RocketConfig.fir@100954.4]
  assign sourceA_io_req_bits_set = _T_602[174:165]; // @[Scheduler.scala 133:18:chipyard.TestHarness.RocketConfig.fir@100954.4]
  assign sourceA_io_req_bits_param = _T_602[164:162]; // @[Scheduler.scala 133:18:chipyard.TestHarness.RocketConfig.fir@100954.4]
  assign sourceA_io_req_bits_source = {_T_253,_T_260}; // @[Scheduler.scala 133:18:chipyard.TestHarness.RocketConfig.fir@100954.4]
  assign sourceA_io_req_bits_block = _T_602[158]; // @[Scheduler.scala 133:18:chipyard.TestHarness.RocketConfig.fir@100954.4]
  assign sourceA_io_a_ready = io_out_a_ready; // @[Scheduler.scala 45:12:chipyard.TestHarness.RocketConfig.fir@100053.4]
  assign sourceB_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100035.4]
  assign sourceB_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100036.4]
  assign sourceB_io_req_valid = _T_602[157]; // @[Scheduler.scala 134:18:chipyard.TestHarness.RocketConfig.fir@100955.4]
  assign sourceB_io_req_bits_param = _T_602[156:154]; // @[Scheduler.scala 134:18:chipyard.TestHarness.RocketConfig.fir@100955.4]
  assign sourceB_io_req_bits_tag = _T_602[153:142]; // @[Scheduler.scala 134:18:chipyard.TestHarness.RocketConfig.fir@100955.4]
  assign sourceB_io_req_bits_set = _T_602[141:132]; // @[Scheduler.scala 134:18:chipyard.TestHarness.RocketConfig.fir@100955.4]
  assign sourceB_io_req_bits_clients = _T_602[131]; // @[Scheduler.scala 134:18:chipyard.TestHarness.RocketConfig.fir@100955.4]
  assign sourceB_io_b_ready = io_in_b_ready; // @[Scheduler.scala 48:11:chipyard.TestHarness.RocketConfig.fir@100056.4]
  assign sourceC_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100039.4]
  assign sourceC_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100040.4]
  assign sourceC_io_req_valid = _T_602[130]; // @[Scheduler.scala 135:18:chipyard.TestHarness.RocketConfig.fir@100956.4]
  assign sourceC_io_req_bits_opcode = _T_602[129:127]; // @[Scheduler.scala 135:18:chipyard.TestHarness.RocketConfig.fir@100956.4]
  assign sourceC_io_req_bits_param = _T_602[126:124]; // @[Scheduler.scala 135:18:chipyard.TestHarness.RocketConfig.fir@100956.4]
  assign sourceC_io_req_bits_source = schedule_c_bits_opcode[1] ? mshr_select : 3'h0; // @[Scheduler.scala 135:18:chipyard.TestHarness.RocketConfig.fir@100956.4]
  assign sourceC_io_req_bits_tag = _T_602[120:109]; // @[Scheduler.scala 135:18:chipyard.TestHarness.RocketConfig.fir@100956.4]
  assign sourceC_io_req_bits_set = _T_602[108:99]; // @[Scheduler.scala 135:18:chipyard.TestHarness.RocketConfig.fir@100956.4]
  assign sourceC_io_req_bits_way = _T_602[98:96]; // @[Scheduler.scala 135:18:chipyard.TestHarness.RocketConfig.fir@100956.4]
  assign sourceC_io_req_bits_dirty = _T_602[95]; // @[Scheduler.scala 135:18:chipyard.TestHarness.RocketConfig.fir@100956.4]
  assign sourceC_io_c_ready = io_out_c_ready; // @[Scheduler.scala 46:12:chipyard.TestHarness.RocketConfig.fir@100054.4]
  assign sourceC_io_bs_adr_ready = bankedStore_io_sourceC_adr_ready; // @[Scheduler.scala 322:30:chipyard.TestHarness.RocketConfig.fir@101735.4]
  assign sourceC_io_bs_dat_data = bankedStore_io_sourceC_dat_data; // @[Scheduler.scala 326:21:chipyard.TestHarness.RocketConfig.fir@101739.4]
  assign sourceC_io_evict_safe = sourceD_io_evict_safe; // @[Scheduler.scala 332:25:chipyard.TestHarness.RocketConfig.fir@101743.4]
  assign sourceD_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100043.4]
  assign sourceD_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100044.4]
  assign sourceD_io_req_valid = _T_602[94]; // @[Scheduler.scala 136:18:chipyard.TestHarness.RocketConfig.fir@100957.4]
  assign sourceD_io_req_bits_prio_0 = _T_602[91]; // @[Scheduler.scala 136:18:chipyard.TestHarness.RocketConfig.fir@100957.4]
  assign sourceD_io_req_bits_prio_2 = _T_602[93]; // @[Scheduler.scala 136:18:chipyard.TestHarness.RocketConfig.fir@100957.4]
  assign sourceD_io_req_bits_opcode = _T_602[89:87]; // @[Scheduler.scala 136:18:chipyard.TestHarness.RocketConfig.fir@100957.4]
  assign sourceD_io_req_bits_param = _T_602[86:84]; // @[Scheduler.scala 136:18:chipyard.TestHarness.RocketConfig.fir@100957.4]
  assign sourceD_io_req_bits_size = _T_602[83:81]; // @[Scheduler.scala 136:18:chipyard.TestHarness.RocketConfig.fir@100957.4]
  assign sourceD_io_req_bits_source = _T_602[80:78]; // @[Scheduler.scala 136:18:chipyard.TestHarness.RocketConfig.fir@100957.4]
  assign sourceD_io_req_bits_offset = _T_602[65:60]; // @[Scheduler.scala 136:18:chipyard.TestHarness.RocketConfig.fir@100957.4]
  assign sourceD_io_req_bits_put = _T_602[59:54]; // @[Scheduler.scala 136:18:chipyard.TestHarness.RocketConfig.fir@100957.4]
  assign sourceD_io_req_bits_set = _T_602[53:44]; // @[Scheduler.scala 136:18:chipyard.TestHarness.RocketConfig.fir@100957.4]
  assign sourceD_io_req_bits_sink = {_T_253,_T_260}; // @[Scheduler.scala 136:18:chipyard.TestHarness.RocketConfig.fir@100957.4]
  assign sourceD_io_req_bits_way = _T_602[40:38]; // @[Scheduler.scala 136:18:chipyard.TestHarness.RocketConfig.fir@100957.4]
  assign sourceD_io_req_bits_bad = _T_602[37]; // @[Scheduler.scala 136:18:chipyard.TestHarness.RocketConfig.fir@100957.4]
  assign sourceD_io_d_ready = io_in_d_ready; // @[Scheduler.scala 49:11:chipyard.TestHarness.RocketConfig.fir@100057.4]
  assign sourceD_io_pb_pop_ready = sinkA_io_pb_pop_ready; // @[Scheduler.scala 312:19:chipyard.TestHarness.RocketConfig.fir@101727.4]
  assign sourceD_io_pb_beat_data = sinkA_io_pb_beat_data; // @[Scheduler.scala 313:22:chipyard.TestHarness.RocketConfig.fir@101728.4]
  assign sourceD_io_pb_beat_mask = sinkA_io_pb_beat_mask; // @[Scheduler.scala 313:22:chipyard.TestHarness.RocketConfig.fir@101728.4]
  assign sourceD_io_pb_beat_corrupt = sinkA_io_pb_beat_corrupt; // @[Scheduler.scala 313:22:chipyard.TestHarness.RocketConfig.fir@101728.4]
  assign sourceD_io_rel_pop_ready = sinkC_io_rel_pop_ready; // @[Scheduler.scala 314:20:chipyard.TestHarness.RocketConfig.fir@101729.4]
  assign sourceD_io_rel_beat_data = sinkC_io_rel_beat_data; // @[Scheduler.scala 315:23:chipyard.TestHarness.RocketConfig.fir@101730.4]
  assign sourceD_io_rel_beat_corrupt = sinkC_io_rel_beat_corrupt; // @[Scheduler.scala 315:23:chipyard.TestHarness.RocketConfig.fir@101730.4]
  assign sourceD_io_bs_radr_ready = bankedStore_io_sourceD_radr_ready; // @[Scheduler.scala 323:31:chipyard.TestHarness.RocketConfig.fir@101736.4]
  assign sourceD_io_bs_rdat_data = bankedStore_io_sourceD_rdat_data; // @[Scheduler.scala 327:22:chipyard.TestHarness.RocketConfig.fir@101740.4]
  assign sourceD_io_bs_wadr_ready = bankedStore_io_sourceD_wadr_ready; // @[Scheduler.scala 324:31:chipyard.TestHarness.RocketConfig.fir@101737.4]
  assign sourceD_io_evict_req_set = sourceC_io_evict_req_set; // @[Scheduler.scala 330:24:chipyard.TestHarness.RocketConfig.fir@101741.4]
  assign sourceD_io_evict_req_way = sourceC_io_evict_req_way; // @[Scheduler.scala 330:24:chipyard.TestHarness.RocketConfig.fir@101741.4]
  assign sourceD_io_grant_req_set = sinkD_io_grant_req_set; // @[Scheduler.scala 331:24:chipyard.TestHarness.RocketConfig.fir@101742.4]
  assign sourceD_io_grant_req_way = sinkD_io_grant_req_way; // @[Scheduler.scala 331:24:chipyard.TestHarness.RocketConfig.fir@101742.4]
  assign sourceE_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100047.4]
  assign sourceE_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100048.4]
  assign sourceE_io_req_valid = _T_602[36]; // @[Scheduler.scala 137:18:chipyard.TestHarness.RocketConfig.fir@100958.4]
  assign sourceE_io_req_bits_sink = _T_602[35:33]; // @[Scheduler.scala 137:18:chipyard.TestHarness.RocketConfig.fir@100958.4]
  assign sourceX_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100051.4]
  assign sourceX_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100052.4]
  assign sourceX_io_req_valid = _T_602[32]; // @[Scheduler.scala 138:18:chipyard.TestHarness.RocketConfig.fir@100959.4]
  assign sourceX_io_x_ready = io_resp_ready; // @[Scheduler.scala 50:11:chipyard.TestHarness.RocketConfig.fir@100058.4]
  assign sinkA_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100061.4]
  assign sinkA_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100062.4]
  assign sinkA_io_req_ready = _T_721 & _T_725; // @[Scheduler.scala 158:22:chipyard.TestHarness.RocketConfig.fir@101000.4]
  assign sinkA_io_a_valid = io_in_a_valid; // @[Scheduler.scala 58:14:chipyard.TestHarness.RocketConfig.fir@100079.4]
  assign sinkA_io_a_bits_opcode = io_in_a_bits_opcode; // @[Scheduler.scala 58:14:chipyard.TestHarness.RocketConfig.fir@100079.4]
  assign sinkA_io_a_bits_param = io_in_a_bits_param; // @[Scheduler.scala 58:14:chipyard.TestHarness.RocketConfig.fir@100079.4]
  assign sinkA_io_a_bits_size = io_in_a_bits_size; // @[Scheduler.scala 58:14:chipyard.TestHarness.RocketConfig.fir@100079.4]
  assign sinkA_io_a_bits_source = io_in_a_bits_source; // @[Scheduler.scala 58:14:chipyard.TestHarness.RocketConfig.fir@100079.4]
  assign sinkA_io_a_bits_address = io_in_a_bits_address; // @[Scheduler.scala 58:14:chipyard.TestHarness.RocketConfig.fir@100079.4]
  assign sinkA_io_a_bits_mask = io_in_a_bits_mask; // @[Scheduler.scala 58:14:chipyard.TestHarness.RocketConfig.fir@100079.4]
  assign sinkA_io_a_bits_data = io_in_a_bits_data; // @[Scheduler.scala 58:14:chipyard.TestHarness.RocketConfig.fir@100079.4]
  assign sinkA_io_a_bits_corrupt = io_in_a_bits_corrupt; // @[Scheduler.scala 58:14:chipyard.TestHarness.RocketConfig.fir@100079.4]
  assign sinkA_io_pb_pop_valid = sourceD_io_pb_pop_valid; // @[Scheduler.scala 312:19:chipyard.TestHarness.RocketConfig.fir@101727.4]
  assign sinkA_io_pb_pop_bits_index = sourceD_io_pb_pop_bits_index; // @[Scheduler.scala 312:19:chipyard.TestHarness.RocketConfig.fir@101727.4]
  assign sinkA_io_pb_pop_bits_last = sourceD_io_pb_pop_bits_last; // @[Scheduler.scala 312:19:chipyard.TestHarness.RocketConfig.fir@101727.4]
  assign sinkC_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100065.4]
  assign sinkC_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100066.4]
  assign sinkC_io_req_ready = directory_io_ready & request_ready; // @[Scheduler.scala 156:22:chipyard.TestHarness.RocketConfig.fir@100990.4]
  assign sinkC_io_c_valid = io_in_c_valid; // @[Scheduler.scala 59:14:chipyard.TestHarness.RocketConfig.fir@100080.4]
  assign sinkC_io_c_bits_opcode = io_in_c_bits_opcode; // @[Scheduler.scala 59:14:chipyard.TestHarness.RocketConfig.fir@100080.4]
  assign sinkC_io_c_bits_param = io_in_c_bits_param; // @[Scheduler.scala 59:14:chipyard.TestHarness.RocketConfig.fir@100080.4]
  assign sinkC_io_c_bits_size = io_in_c_bits_size; // @[Scheduler.scala 59:14:chipyard.TestHarness.RocketConfig.fir@100080.4]
  assign sinkC_io_c_bits_source = io_in_c_bits_source; // @[Scheduler.scala 59:14:chipyard.TestHarness.RocketConfig.fir@100080.4]
  assign sinkC_io_c_bits_address = io_in_c_bits_address; // @[Scheduler.scala 59:14:chipyard.TestHarness.RocketConfig.fir@100080.4]
  assign sinkC_io_c_bits_data = io_in_c_bits_data; // @[Scheduler.scala 59:14:chipyard.TestHarness.RocketConfig.fir@100080.4]
  assign sinkC_io_c_bits_corrupt = io_in_c_bits_corrupt; // @[Scheduler.scala 59:14:chipyard.TestHarness.RocketConfig.fir@100080.4]
  assign sinkC_io_way = _T_1238 ? bc_mshr_io_status_bits_way : _T_1257; // @[Scheduler.scala 303:16:chipyard.TestHarness.RocketConfig.fir@101706.4]
  assign sinkC_io_bs_adr_ready = bankedStore_io_sinkC_adr_ready; // @[Scheduler.scala 318:28:chipyard.TestHarness.RocketConfig.fir@101731.4]
  assign sinkC_io_rel_pop_valid = sourceD_io_rel_pop_valid; // @[Scheduler.scala 314:20:chipyard.TestHarness.RocketConfig.fir@101729.4]
  assign sinkC_io_rel_pop_bits_index = sourceD_io_rel_pop_bits_index; // @[Scheduler.scala 314:20:chipyard.TestHarness.RocketConfig.fir@101729.4]
  assign sinkC_io_rel_pop_bits_last = sourceD_io_rel_pop_bits_last; // @[Scheduler.scala 314:20:chipyard.TestHarness.RocketConfig.fir@101729.4]
  assign sinkD_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100069.4]
  assign sinkD_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100070.4]
  assign sinkD_io_d_valid = io_out_d_valid; // @[Scheduler.scala 61:14:chipyard.TestHarness.RocketConfig.fir@100082.4]
  assign sinkD_io_d_bits_opcode = io_out_d_bits_opcode; // @[Scheduler.scala 61:14:chipyard.TestHarness.RocketConfig.fir@100082.4]
  assign sinkD_io_d_bits_param = io_out_d_bits_param; // @[Scheduler.scala 61:14:chipyard.TestHarness.RocketConfig.fir@100082.4]
  assign sinkD_io_d_bits_size = io_out_d_bits_size; // @[Scheduler.scala 61:14:chipyard.TestHarness.RocketConfig.fir@100082.4]
  assign sinkD_io_d_bits_source = io_out_d_bits_source; // @[Scheduler.scala 61:14:chipyard.TestHarness.RocketConfig.fir@100082.4]
  assign sinkD_io_d_bits_sink = io_out_d_bits_sink; // @[Scheduler.scala 61:14:chipyard.TestHarness.RocketConfig.fir@100082.4]
  assign sinkD_io_d_bits_denied = io_out_d_bits_denied; // @[Scheduler.scala 61:14:chipyard.TestHarness.RocketConfig.fir@100082.4]
  assign sinkD_io_d_bits_data = io_out_d_bits_data; // @[Scheduler.scala 61:14:chipyard.TestHarness.RocketConfig.fir@100082.4]
  assign sinkD_io_d_bits_corrupt = io_out_d_bits_corrupt; // @[Scheduler.scala 61:14:chipyard.TestHarness.RocketConfig.fir@100082.4]
  assign sinkD_io_way = 3'h6 == sinkD_io_source ? _T_1260_6 : _GEN_132; // @[Scheduler.scala 308:16:chipyard.TestHarness.RocketConfig.fir@101716.4]
  assign sinkD_io_set = 3'h6 == sinkD_io_source ? _T_1261_6 : _GEN_139; // @[Scheduler.scala 309:16:chipyard.TestHarness.RocketConfig.fir@101726.4]
  assign sinkD_io_bs_adr_ready = bankedStore_io_sinkD_adr_ready; // @[Scheduler.scala 320:28:chipyard.TestHarness.RocketConfig.fir@101733.4]
  assign sinkD_io_grant_safe = sourceD_io_grant_safe; // @[Scheduler.scala 333:25:chipyard.TestHarness.RocketConfig.fir@101744.4]
  assign sinkE_io_e_valid = io_in_e_valid; // @[Scheduler.scala 60:14:chipyard.TestHarness.RocketConfig.fir@100081.4]
  assign sinkE_io_e_bits_sink = io_in_e_bits_sink; // @[Scheduler.scala 60:14:chipyard.TestHarness.RocketConfig.fir@100081.4]
  assign sinkX_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100077.4]
  assign sinkX_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100078.4]
  assign sinkX_io_req_ready = _T_718 & _T_720; // @[Scheduler.scala 157:22:chipyard.TestHarness.RocketConfig.fir@100994.4]
  assign sinkX_io_x_valid = io_req_valid; // @[Scheduler.scala 62:14:chipyard.TestHarness.RocketConfig.fir@100083.4]
  assign sinkX_io_x_bits_address = io_req_bits_address; // @[Scheduler.scala 62:14:chipyard.TestHarness.RocketConfig.fir@100083.4]
  assign directory_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100087.4]
  assign directory_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100088.4]
  assign directory_io_write_valid = _T_602[30]; // @[Scheduler.scala 139:22:chipyard.TestHarness.RocketConfig.fir@100960.4]
  assign directory_io_write_bits_set = _T_602[29:20]; // @[Scheduler.scala 139:22:chipyard.TestHarness.RocketConfig.fir@100960.4]
  assign directory_io_write_bits_way = _T_602[19:17]; // @[Scheduler.scala 139:22:chipyard.TestHarness.RocketConfig.fir@100960.4]
  assign directory_io_write_bits_data_dirty = _T_602[16]; // @[Scheduler.scala 139:22:chipyard.TestHarness.RocketConfig.fir@100960.4]
  assign directory_io_write_bits_data_state = _T_602[15:14]; // @[Scheduler.scala 139:22:chipyard.TestHarness.RocketConfig.fir@100960.4]
  assign directory_io_write_bits_data_clients = _T_602[13]; // @[Scheduler.scala 139:22:chipyard.TestHarness.RocketConfig.fir@100960.4]
  assign directory_io_write_bits_data_tag = _T_602[12:1]; // @[Scheduler.scala 139:22:chipyard.TestHarness.RocketConfig.fir@100960.4]
  assign directory_io_read_valid = mshr_uses_directory | alloc_uses_directory; // @[Scheduler.scala 254:27:chipyard.TestHarness.RocketConfig.fir@101450.4]
  assign directory_io_read_bits_set = mshr_uses_directory_for_lb ? scheduleSet : request_bits_set; // @[Scheduler.scala 255:30:chipyard.TestHarness.RocketConfig.fir@101452.4]
  assign directory_io_read_bits_tag = mshr_uses_directory_for_lb ? requests_io_data_tag : request_bits_tag; // @[Scheduler.scala 256:30:chipyard.TestHarness.RocketConfig.fir@101454.4]
  assign bankedStore_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100091.4]
  assign bankedStore_io_sinkC_adr_valid = sinkC_io_bs_adr_valid; // @[Scheduler.scala 318:28:chipyard.TestHarness.RocketConfig.fir@101731.4]
  assign bankedStore_io_sinkC_adr_bits_noop = sinkC_io_bs_adr_bits_noop; // @[Scheduler.scala 318:28:chipyard.TestHarness.RocketConfig.fir@101731.4]
  assign bankedStore_io_sinkC_adr_bits_way = sinkC_io_bs_adr_bits_way; // @[Scheduler.scala 318:28:chipyard.TestHarness.RocketConfig.fir@101731.4]
  assign bankedStore_io_sinkC_adr_bits_set = sinkC_io_bs_adr_bits_set; // @[Scheduler.scala 318:28:chipyard.TestHarness.RocketConfig.fir@101731.4]
  assign bankedStore_io_sinkC_adr_bits_beat = sinkC_io_bs_adr_bits_beat; // @[Scheduler.scala 318:28:chipyard.TestHarness.RocketConfig.fir@101731.4]
  assign bankedStore_io_sinkC_adr_bits_mask = sinkC_io_bs_adr_bits_mask; // @[Scheduler.scala 318:28:chipyard.TestHarness.RocketConfig.fir@101731.4]
  assign bankedStore_io_sinkC_dat_data = sinkC_io_bs_dat_data; // @[Scheduler.scala 319:28:chipyard.TestHarness.RocketConfig.fir@101732.4]
  assign bankedStore_io_sinkD_adr_valid = sinkD_io_bs_adr_valid; // @[Scheduler.scala 320:28:chipyard.TestHarness.RocketConfig.fir@101733.4]
  assign bankedStore_io_sinkD_adr_bits_noop = sinkD_io_bs_adr_bits_noop; // @[Scheduler.scala 320:28:chipyard.TestHarness.RocketConfig.fir@101733.4]
  assign bankedStore_io_sinkD_adr_bits_way = sinkD_io_bs_adr_bits_way; // @[Scheduler.scala 320:28:chipyard.TestHarness.RocketConfig.fir@101733.4]
  assign bankedStore_io_sinkD_adr_bits_set = sinkD_io_bs_adr_bits_set; // @[Scheduler.scala 320:28:chipyard.TestHarness.RocketConfig.fir@101733.4]
  assign bankedStore_io_sinkD_adr_bits_beat = sinkD_io_bs_adr_bits_beat; // @[Scheduler.scala 320:28:chipyard.TestHarness.RocketConfig.fir@101733.4]
  assign bankedStore_io_sinkD_dat_data = sinkD_io_bs_dat_data; // @[Scheduler.scala 321:28:chipyard.TestHarness.RocketConfig.fir@101734.4]
  assign bankedStore_io_sourceC_adr_valid = sourceC_io_bs_adr_valid; // @[Scheduler.scala 322:30:chipyard.TestHarness.RocketConfig.fir@101735.4]
  assign bankedStore_io_sourceC_adr_bits_way = sourceC_io_bs_adr_bits_way; // @[Scheduler.scala 322:30:chipyard.TestHarness.RocketConfig.fir@101735.4]
  assign bankedStore_io_sourceC_adr_bits_set = sourceC_io_bs_adr_bits_set; // @[Scheduler.scala 322:30:chipyard.TestHarness.RocketConfig.fir@101735.4]
  assign bankedStore_io_sourceC_adr_bits_beat = sourceC_io_bs_adr_bits_beat; // @[Scheduler.scala 322:30:chipyard.TestHarness.RocketConfig.fir@101735.4]
  assign bankedStore_io_sourceD_radr_valid = sourceD_io_bs_radr_valid; // @[Scheduler.scala 323:31:chipyard.TestHarness.RocketConfig.fir@101736.4]
  assign bankedStore_io_sourceD_radr_bits_way = sourceD_io_bs_radr_bits_way; // @[Scheduler.scala 323:31:chipyard.TestHarness.RocketConfig.fir@101736.4]
  assign bankedStore_io_sourceD_radr_bits_set = sourceD_io_bs_radr_bits_set; // @[Scheduler.scala 323:31:chipyard.TestHarness.RocketConfig.fir@101736.4]
  assign bankedStore_io_sourceD_radr_bits_beat = sourceD_io_bs_radr_bits_beat; // @[Scheduler.scala 323:31:chipyard.TestHarness.RocketConfig.fir@101736.4]
  assign bankedStore_io_sourceD_radr_bits_mask = sourceD_io_bs_radr_bits_mask; // @[Scheduler.scala 323:31:chipyard.TestHarness.RocketConfig.fir@101736.4]
  assign bankedStore_io_sourceD_wadr_valid = sourceD_io_bs_wadr_valid; // @[Scheduler.scala 324:31:chipyard.TestHarness.RocketConfig.fir@101737.4]
  assign bankedStore_io_sourceD_wadr_bits_way = sourceD_io_bs_wadr_bits_way; // @[Scheduler.scala 324:31:chipyard.TestHarness.RocketConfig.fir@101737.4]
  assign bankedStore_io_sourceD_wadr_bits_set = sourceD_io_bs_wadr_bits_set; // @[Scheduler.scala 324:31:chipyard.TestHarness.RocketConfig.fir@101737.4]
  assign bankedStore_io_sourceD_wadr_bits_beat = sourceD_io_bs_wadr_bits_beat; // @[Scheduler.scala 324:31:chipyard.TestHarness.RocketConfig.fir@101737.4]
  assign bankedStore_io_sourceD_wadr_bits_mask = sourceD_io_bs_wadr_bits_mask; // @[Scheduler.scala 324:31:chipyard.TestHarness.RocketConfig.fir@101737.4]
  assign bankedStore_io_sourceD_wdat_data = sourceD_io_bs_wdat_data; // @[Scheduler.scala 325:31:chipyard.TestHarness.RocketConfig.fir@101738.4]
  assign requests_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100095.4]
  assign requests_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100096.4]
  assign requests_io_push_valid = _T_844 & _T_1093; // @[Scheduler.scala 259:26:chipyard.TestHarness.RocketConfig.fir@101458.4]
  assign requests_io_push_bits_index = _GEN_152 | _T_1148; // @[Scheduler.scala 261:31:chipyard.TestHarness.RocketConfig.fir@101518.4]
  assign requests_io_push_bits_data_prio_0 = sinkC_io_req_valid ? 1'h0 : 1'h1; // @[Scheduler.scala 260:31:chipyard.TestHarness.RocketConfig.fir@101459.4]
  assign requests_io_push_bits_data_prio_2 = sinkC_io_req_valid; // @[Scheduler.scala 260:31:chipyard.TestHarness.RocketConfig.fir@101459.4]
  assign requests_io_push_bits_data_control = sinkC_io_req_valid ? 1'h0 : _T_716_control; // @[Scheduler.scala 260:31:chipyard.TestHarness.RocketConfig.fir@101459.4]
  assign requests_io_push_bits_data_opcode = sinkC_io_req_valid ? sinkC_io_req_bits_opcode : _T_716_opcode; // @[Scheduler.scala 260:31:chipyard.TestHarness.RocketConfig.fir@101459.4]
  assign requests_io_push_bits_data_param = sinkC_io_req_valid ? sinkC_io_req_bits_param : _T_716_param; // @[Scheduler.scala 260:31:chipyard.TestHarness.RocketConfig.fir@101459.4]
  assign requests_io_push_bits_data_size = sinkC_io_req_valid ? sinkC_io_req_bits_size : _T_716_size; // @[Scheduler.scala 260:31:chipyard.TestHarness.RocketConfig.fir@101459.4]
  assign requests_io_push_bits_data_source = sinkC_io_req_valid ? sinkC_io_req_bits_source : _T_716_source; // @[Scheduler.scala 260:31:chipyard.TestHarness.RocketConfig.fir@101459.4]
  assign requests_io_push_bits_data_tag = sinkC_io_req_valid ? sinkC_io_req_bits_tag : _T_716_tag; // @[Scheduler.scala 260:31:chipyard.TestHarness.RocketConfig.fir@101459.4]
  assign requests_io_push_bits_data_offset = sinkC_io_req_valid ? sinkC_io_req_bits_offset : _T_716_offset; // @[Scheduler.scala 260:31:chipyard.TestHarness.RocketConfig.fir@101459.4]
  assign requests_io_push_bits_data_put = sinkC_io_req_valid ? sinkC_io_req_bits_put : _T_716_put; // @[Scheduler.scala 260:31:chipyard.TestHarness.RocketConfig.fir@101459.4]
  assign requests_io_pop_valid = _T_1062 & _T_866; // @[Scheduler.scala 231:25:chipyard.TestHarness.RocketConfig.fir@101410.4]
  assign requests_io_pop_bits = {_T_1044,_T_1061}; // @[Scheduler.scala 232:25:chipyard.TestHarness.RocketConfig.fir@101411.4]
  assign abc_mshrs_0_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100099.4]
  assign abc_mshrs_0_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100100.4]
  assign abc_mshrs_0_io_allocate_valid = _T_1178 | _T_895; // @[Scheduler.scala 225:25:chipyard.TestHarness.RocketConfig.fir@101199.4 Scheduler.scala 270:27:chipyard.TestHarness.RocketConfig.fir@101548.6]
  assign abc_mshrs_0_io_allocate_bits_prio_0 = _T_1178 ? request_bits_prio_0 : _T_893_prio_0; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101194.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101549.6]
  assign abc_mshrs_0_io_allocate_bits_prio_1 = _T_1178 ? 1'h0 : _T_893_prio_1; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101194.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101549.6]
  assign abc_mshrs_0_io_allocate_bits_prio_2 = _T_1178 ? request_bits_prio_2 : _T_893_prio_2; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101194.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101549.6]
  assign abc_mshrs_0_io_allocate_bits_control = _T_1178 ? request_bits_control : _T_893_control; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101194.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101549.6]
  assign abc_mshrs_0_io_allocate_bits_opcode = _T_1178 ? request_bits_opcode : _T_893_opcode; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101194.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101549.6]
  assign abc_mshrs_0_io_allocate_bits_param = _T_1178 ? request_bits_param : _T_893_param; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101194.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101549.6]
  assign abc_mshrs_0_io_allocate_bits_size = _T_1178 ? request_bits_size : _T_893_size; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101194.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101549.6]
  assign abc_mshrs_0_io_allocate_bits_source = _T_1178 ? request_bits_source : _T_893_source; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101194.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101549.6]
  assign abc_mshrs_0_io_allocate_bits_tag = _T_1178 ? request_bits_tag : _T_893_tag; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101194.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101549.6]
  assign abc_mshrs_0_io_allocate_bits_offset = _T_1178 ? request_bits_offset : _T_893_offset; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101194.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101549.6]
  assign abc_mshrs_0_io_allocate_bits_put = _T_1178 ? request_bits_put : _T_893_put; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101194.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101549.6]
  assign abc_mshrs_0_io_allocate_bits_set = _T_1178 ? request_bits_set : abc_mshrs_0_io_status_bits_set; // @[Scheduler.scala 223:28:chipyard.TestHarness.RocketConfig.fir@101195.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101549.6]
  assign abc_mshrs_0_io_allocate_bits_repeat = _T_1178 ? 1'h0 : _T_894; // @[Scheduler.scala 224:31:chipyard.TestHarness.RocketConfig.fir@101197.4 Scheduler.scala 272:33:chipyard.TestHarness.RocketConfig.fir@101550.6]
  assign abc_mshrs_0_io_directory_valid = directoryFanout[0]; // @[Scheduler.scala 298:26:chipyard.TestHarness.RocketConfig.fir@101662.4]
  assign abc_mshrs_0_io_directory_bits_dirty = directory_io_result_bits_dirty; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101663.4]
  assign abc_mshrs_0_io_directory_bits_state = directory_io_result_bits_state; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101663.4]
  assign abc_mshrs_0_io_directory_bits_clients = directory_io_result_bits_clients; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101663.4]
  assign abc_mshrs_0_io_directory_bits_tag = directory_io_result_bits_tag; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101663.4]
  assign abc_mshrs_0_io_directory_bits_hit = directory_io_result_bits_hit; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101663.4]
  assign abc_mshrs_0_io_directory_bits_way = directory_io_result_bits_way; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101663.4]
  assign abc_mshrs_0_io_schedule_ready = mshr_selectOH[0]; // @[Scheduler.scala 213:25:chipyard.TestHarness.RocketConfig.fir@101171.4]
  assign abc_mshrs_0_io_sinkc_valid = sinkC_io_resp_valid & _T; // @[Scheduler.scala 77:22:chipyard.TestHarness.RocketConfig.fir@100129.4]
  assign abc_mshrs_0_io_sinkc_bits_last = sinkC_io_resp_bits_last; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100136.4]
  assign abc_mshrs_0_io_sinkc_bits_tag = sinkC_io_resp_bits_tag; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100136.4]
  assign abc_mshrs_0_io_sinkc_bits_source = sinkC_io_resp_bits_source; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100136.4]
  assign abc_mshrs_0_io_sinkc_bits_param = sinkC_io_resp_bits_param; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100136.4]
  assign abc_mshrs_0_io_sinkc_bits_data = sinkC_io_resp_bits_data; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100136.4]
  assign abc_mshrs_0_io_sinkd_valid = sinkD_io_resp_valid & _T_2; // @[Scheduler.scala 78:22:chipyard.TestHarness.RocketConfig.fir@100132.4]
  assign abc_mshrs_0_io_sinkd_bits_last = sinkD_io_resp_bits_last; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100137.4]
  assign abc_mshrs_0_io_sinkd_bits_opcode = sinkD_io_resp_bits_opcode; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100137.4]
  assign abc_mshrs_0_io_sinkd_bits_param = sinkD_io_resp_bits_param; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100137.4]
  assign abc_mshrs_0_io_sinkd_bits_sink = sinkD_io_resp_bits_sink; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100137.4]
  assign abc_mshrs_0_io_sinkd_bits_denied = sinkD_io_resp_bits_denied; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100137.4]
  assign abc_mshrs_0_io_sinke_valid = sinkE_io_resp_valid & _T_4; // @[Scheduler.scala 79:22:chipyard.TestHarness.RocketConfig.fir@100135.4]
  assign abc_mshrs_0_io_nestedwb_set = mshr_selectOH[6] ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100139.4]
  assign abc_mshrs_0_io_nestedwb_tag = mshr_selectOH[6] ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100139.4]
  assign abc_mshrs_0_io_nestedwb_b_toN = _T_704 & _T_705; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100139.4]
  assign abc_mshrs_0_io_nestedwb_b_toB = _T_704 & _T_708; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100139.4]
  assign abc_mshrs_0_io_nestedwb_b_clr_dirty = mshr_selectOH[5] & bc_mshr_io_schedule_bits_dir_valid; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100139.4]
  assign abc_mshrs_0_io_nestedwb_c_set_dirty = _T_711 & c_mshr_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100139.4]
  assign abc_mshrs_1_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100103.4]
  assign abc_mshrs_1_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100104.4]
  assign abc_mshrs_1_io_allocate_valid = _T_1182 | _T_918; // @[Scheduler.scala 225:25:chipyard.TestHarness.RocketConfig.fir@101229.4 Scheduler.scala 270:27:chipyard.TestHarness.RocketConfig.fir@101557.6]
  assign abc_mshrs_1_io_allocate_bits_prio_0 = _T_1182 ? request_bits_prio_0 : _T_916_prio_0; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101224.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101558.6]
  assign abc_mshrs_1_io_allocate_bits_prio_1 = _T_1182 ? 1'h0 : _T_916_prio_1; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101224.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101558.6]
  assign abc_mshrs_1_io_allocate_bits_prio_2 = _T_1182 ? request_bits_prio_2 : _T_916_prio_2; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101224.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101558.6]
  assign abc_mshrs_1_io_allocate_bits_control = _T_1182 ? request_bits_control : _T_916_control; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101224.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101558.6]
  assign abc_mshrs_1_io_allocate_bits_opcode = _T_1182 ? request_bits_opcode : _T_916_opcode; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101224.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101558.6]
  assign abc_mshrs_1_io_allocate_bits_param = _T_1182 ? request_bits_param : _T_916_param; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101224.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101558.6]
  assign abc_mshrs_1_io_allocate_bits_size = _T_1182 ? request_bits_size : _T_916_size; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101224.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101558.6]
  assign abc_mshrs_1_io_allocate_bits_source = _T_1182 ? request_bits_source : _T_916_source; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101224.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101558.6]
  assign abc_mshrs_1_io_allocate_bits_tag = _T_1182 ? request_bits_tag : _T_916_tag; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101224.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101558.6]
  assign abc_mshrs_1_io_allocate_bits_offset = _T_1182 ? request_bits_offset : _T_916_offset; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101224.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101558.6]
  assign abc_mshrs_1_io_allocate_bits_put = _T_1182 ? request_bits_put : _T_916_put; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101224.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101558.6]
  assign abc_mshrs_1_io_allocate_bits_set = _T_1182 ? request_bits_set : abc_mshrs_1_io_status_bits_set; // @[Scheduler.scala 223:28:chipyard.TestHarness.RocketConfig.fir@101225.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101558.6]
  assign abc_mshrs_1_io_allocate_bits_repeat = _T_1182 ? 1'h0 : _T_917; // @[Scheduler.scala 224:31:chipyard.TestHarness.RocketConfig.fir@101227.4 Scheduler.scala 272:33:chipyard.TestHarness.RocketConfig.fir@101559.6]
  assign abc_mshrs_1_io_directory_valid = directoryFanout[1]; // @[Scheduler.scala 298:26:chipyard.TestHarness.RocketConfig.fir@101665.4]
  assign abc_mshrs_1_io_directory_bits_dirty = directory_io_result_bits_dirty; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101666.4]
  assign abc_mshrs_1_io_directory_bits_state = directory_io_result_bits_state; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101666.4]
  assign abc_mshrs_1_io_directory_bits_clients = directory_io_result_bits_clients; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101666.4]
  assign abc_mshrs_1_io_directory_bits_tag = directory_io_result_bits_tag; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101666.4]
  assign abc_mshrs_1_io_directory_bits_hit = directory_io_result_bits_hit; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101666.4]
  assign abc_mshrs_1_io_directory_bits_way = directory_io_result_bits_way; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101666.4]
  assign abc_mshrs_1_io_schedule_ready = mshr_selectOH[1]; // @[Scheduler.scala 213:25:chipyard.TestHarness.RocketConfig.fir@101201.4]
  assign abc_mshrs_1_io_sinkc_valid = sinkC_io_resp_valid & _T_6; // @[Scheduler.scala 77:22:chipyard.TestHarness.RocketConfig.fir@100142.4]
  assign abc_mshrs_1_io_sinkc_bits_last = sinkC_io_resp_bits_last; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100149.4]
  assign abc_mshrs_1_io_sinkc_bits_tag = sinkC_io_resp_bits_tag; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100149.4]
  assign abc_mshrs_1_io_sinkc_bits_source = sinkC_io_resp_bits_source; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100149.4]
  assign abc_mshrs_1_io_sinkc_bits_param = sinkC_io_resp_bits_param; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100149.4]
  assign abc_mshrs_1_io_sinkc_bits_data = sinkC_io_resp_bits_data; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100149.4]
  assign abc_mshrs_1_io_sinkd_valid = sinkD_io_resp_valid & _T_8; // @[Scheduler.scala 78:22:chipyard.TestHarness.RocketConfig.fir@100145.4]
  assign abc_mshrs_1_io_sinkd_bits_last = sinkD_io_resp_bits_last; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100150.4]
  assign abc_mshrs_1_io_sinkd_bits_opcode = sinkD_io_resp_bits_opcode; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100150.4]
  assign abc_mshrs_1_io_sinkd_bits_param = sinkD_io_resp_bits_param; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100150.4]
  assign abc_mshrs_1_io_sinkd_bits_sink = sinkD_io_resp_bits_sink; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100150.4]
  assign abc_mshrs_1_io_sinkd_bits_denied = sinkD_io_resp_bits_denied; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100150.4]
  assign abc_mshrs_1_io_sinke_valid = sinkE_io_resp_valid & _T_10; // @[Scheduler.scala 79:22:chipyard.TestHarness.RocketConfig.fir@100148.4]
  assign abc_mshrs_1_io_nestedwb_set = mshr_selectOH[6] ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100152.4]
  assign abc_mshrs_1_io_nestedwb_tag = mshr_selectOH[6] ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100152.4]
  assign abc_mshrs_1_io_nestedwb_b_toN = _T_704 & _T_705; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100152.4]
  assign abc_mshrs_1_io_nestedwb_b_toB = _T_704 & _T_708; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100152.4]
  assign abc_mshrs_1_io_nestedwb_b_clr_dirty = mshr_selectOH[5] & bc_mshr_io_schedule_bits_dir_valid; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100152.4]
  assign abc_mshrs_1_io_nestedwb_c_set_dirty = _T_711 & c_mshr_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100152.4]
  assign abc_mshrs_2_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100107.4]
  assign abc_mshrs_2_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100108.4]
  assign abc_mshrs_2_io_allocate_valid = _T_1186 | _T_941; // @[Scheduler.scala 225:25:chipyard.TestHarness.RocketConfig.fir@101259.4 Scheduler.scala 270:27:chipyard.TestHarness.RocketConfig.fir@101566.6]
  assign abc_mshrs_2_io_allocate_bits_prio_0 = _T_1186 ? request_bits_prio_0 : _T_939_prio_0; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101254.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101567.6]
  assign abc_mshrs_2_io_allocate_bits_prio_1 = _T_1186 ? 1'h0 : _T_939_prio_1; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101254.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101567.6]
  assign abc_mshrs_2_io_allocate_bits_prio_2 = _T_1186 ? request_bits_prio_2 : _T_939_prio_2; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101254.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101567.6]
  assign abc_mshrs_2_io_allocate_bits_control = _T_1186 ? request_bits_control : _T_939_control; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101254.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101567.6]
  assign abc_mshrs_2_io_allocate_bits_opcode = _T_1186 ? request_bits_opcode : _T_939_opcode; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101254.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101567.6]
  assign abc_mshrs_2_io_allocate_bits_param = _T_1186 ? request_bits_param : _T_939_param; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101254.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101567.6]
  assign abc_mshrs_2_io_allocate_bits_size = _T_1186 ? request_bits_size : _T_939_size; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101254.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101567.6]
  assign abc_mshrs_2_io_allocate_bits_source = _T_1186 ? request_bits_source : _T_939_source; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101254.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101567.6]
  assign abc_mshrs_2_io_allocate_bits_tag = _T_1186 ? request_bits_tag : _T_939_tag; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101254.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101567.6]
  assign abc_mshrs_2_io_allocate_bits_offset = _T_1186 ? request_bits_offset : _T_939_offset; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101254.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101567.6]
  assign abc_mshrs_2_io_allocate_bits_put = _T_1186 ? request_bits_put : _T_939_put; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101254.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101567.6]
  assign abc_mshrs_2_io_allocate_bits_set = _T_1186 ? request_bits_set : abc_mshrs_2_io_status_bits_set; // @[Scheduler.scala 223:28:chipyard.TestHarness.RocketConfig.fir@101255.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101567.6]
  assign abc_mshrs_2_io_allocate_bits_repeat = _T_1186 ? 1'h0 : _T_940; // @[Scheduler.scala 224:31:chipyard.TestHarness.RocketConfig.fir@101257.4 Scheduler.scala 272:33:chipyard.TestHarness.RocketConfig.fir@101568.6]
  assign abc_mshrs_2_io_directory_valid = directoryFanout[2]; // @[Scheduler.scala 298:26:chipyard.TestHarness.RocketConfig.fir@101668.4]
  assign abc_mshrs_2_io_directory_bits_dirty = directory_io_result_bits_dirty; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101669.4]
  assign abc_mshrs_2_io_directory_bits_state = directory_io_result_bits_state; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101669.4]
  assign abc_mshrs_2_io_directory_bits_clients = directory_io_result_bits_clients; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101669.4]
  assign abc_mshrs_2_io_directory_bits_tag = directory_io_result_bits_tag; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101669.4]
  assign abc_mshrs_2_io_directory_bits_hit = directory_io_result_bits_hit; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101669.4]
  assign abc_mshrs_2_io_directory_bits_way = directory_io_result_bits_way; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101669.4]
  assign abc_mshrs_2_io_schedule_ready = mshr_selectOH[2]; // @[Scheduler.scala 213:25:chipyard.TestHarness.RocketConfig.fir@101231.4]
  assign abc_mshrs_2_io_sinkc_valid = sinkC_io_resp_valid & _T_12; // @[Scheduler.scala 77:22:chipyard.TestHarness.RocketConfig.fir@100155.4]
  assign abc_mshrs_2_io_sinkc_bits_last = sinkC_io_resp_bits_last; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100162.4]
  assign abc_mshrs_2_io_sinkc_bits_tag = sinkC_io_resp_bits_tag; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100162.4]
  assign abc_mshrs_2_io_sinkc_bits_source = sinkC_io_resp_bits_source; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100162.4]
  assign abc_mshrs_2_io_sinkc_bits_param = sinkC_io_resp_bits_param; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100162.4]
  assign abc_mshrs_2_io_sinkc_bits_data = sinkC_io_resp_bits_data; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100162.4]
  assign abc_mshrs_2_io_sinkd_valid = sinkD_io_resp_valid & _T_14; // @[Scheduler.scala 78:22:chipyard.TestHarness.RocketConfig.fir@100158.4]
  assign abc_mshrs_2_io_sinkd_bits_last = sinkD_io_resp_bits_last; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100163.4]
  assign abc_mshrs_2_io_sinkd_bits_opcode = sinkD_io_resp_bits_opcode; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100163.4]
  assign abc_mshrs_2_io_sinkd_bits_param = sinkD_io_resp_bits_param; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100163.4]
  assign abc_mshrs_2_io_sinkd_bits_sink = sinkD_io_resp_bits_sink; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100163.4]
  assign abc_mshrs_2_io_sinkd_bits_denied = sinkD_io_resp_bits_denied; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100163.4]
  assign abc_mshrs_2_io_sinke_valid = sinkE_io_resp_valid & _T_16; // @[Scheduler.scala 79:22:chipyard.TestHarness.RocketConfig.fir@100161.4]
  assign abc_mshrs_2_io_nestedwb_set = mshr_selectOH[6] ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100165.4]
  assign abc_mshrs_2_io_nestedwb_tag = mshr_selectOH[6] ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100165.4]
  assign abc_mshrs_2_io_nestedwb_b_toN = _T_704 & _T_705; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100165.4]
  assign abc_mshrs_2_io_nestedwb_b_toB = _T_704 & _T_708; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100165.4]
  assign abc_mshrs_2_io_nestedwb_b_clr_dirty = mshr_selectOH[5] & bc_mshr_io_schedule_bits_dir_valid; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100165.4]
  assign abc_mshrs_2_io_nestedwb_c_set_dirty = _T_711 & c_mshr_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100165.4]
  assign abc_mshrs_3_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100111.4]
  assign abc_mshrs_3_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100112.4]
  assign abc_mshrs_3_io_allocate_valid = _T_1190 | _T_964; // @[Scheduler.scala 225:25:chipyard.TestHarness.RocketConfig.fir@101289.4 Scheduler.scala 270:27:chipyard.TestHarness.RocketConfig.fir@101575.6]
  assign abc_mshrs_3_io_allocate_bits_prio_0 = _T_1190 ? request_bits_prio_0 : _T_962_prio_0; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101284.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101576.6]
  assign abc_mshrs_3_io_allocate_bits_prio_1 = _T_1190 ? 1'h0 : _T_962_prio_1; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101284.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101576.6]
  assign abc_mshrs_3_io_allocate_bits_prio_2 = _T_1190 ? request_bits_prio_2 : _T_962_prio_2; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101284.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101576.6]
  assign abc_mshrs_3_io_allocate_bits_control = _T_1190 ? request_bits_control : _T_962_control; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101284.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101576.6]
  assign abc_mshrs_3_io_allocate_bits_opcode = _T_1190 ? request_bits_opcode : _T_962_opcode; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101284.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101576.6]
  assign abc_mshrs_3_io_allocate_bits_param = _T_1190 ? request_bits_param : _T_962_param; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101284.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101576.6]
  assign abc_mshrs_3_io_allocate_bits_size = _T_1190 ? request_bits_size : _T_962_size; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101284.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101576.6]
  assign abc_mshrs_3_io_allocate_bits_source = _T_1190 ? request_bits_source : _T_962_source; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101284.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101576.6]
  assign abc_mshrs_3_io_allocate_bits_tag = _T_1190 ? request_bits_tag : _T_962_tag; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101284.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101576.6]
  assign abc_mshrs_3_io_allocate_bits_offset = _T_1190 ? request_bits_offset : _T_962_offset; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101284.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101576.6]
  assign abc_mshrs_3_io_allocate_bits_put = _T_1190 ? request_bits_put : _T_962_put; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101284.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101576.6]
  assign abc_mshrs_3_io_allocate_bits_set = _T_1190 ? request_bits_set : abc_mshrs_3_io_status_bits_set; // @[Scheduler.scala 223:28:chipyard.TestHarness.RocketConfig.fir@101285.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101576.6]
  assign abc_mshrs_3_io_allocate_bits_repeat = _T_1190 ? 1'h0 : _T_963; // @[Scheduler.scala 224:31:chipyard.TestHarness.RocketConfig.fir@101287.4 Scheduler.scala 272:33:chipyard.TestHarness.RocketConfig.fir@101577.6]
  assign abc_mshrs_3_io_directory_valid = directoryFanout[3]; // @[Scheduler.scala 298:26:chipyard.TestHarness.RocketConfig.fir@101671.4]
  assign abc_mshrs_3_io_directory_bits_dirty = directory_io_result_bits_dirty; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101672.4]
  assign abc_mshrs_3_io_directory_bits_state = directory_io_result_bits_state; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101672.4]
  assign abc_mshrs_3_io_directory_bits_clients = directory_io_result_bits_clients; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101672.4]
  assign abc_mshrs_3_io_directory_bits_tag = directory_io_result_bits_tag; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101672.4]
  assign abc_mshrs_3_io_directory_bits_hit = directory_io_result_bits_hit; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101672.4]
  assign abc_mshrs_3_io_directory_bits_way = directory_io_result_bits_way; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101672.4]
  assign abc_mshrs_3_io_schedule_ready = mshr_selectOH[3]; // @[Scheduler.scala 213:25:chipyard.TestHarness.RocketConfig.fir@101261.4]
  assign abc_mshrs_3_io_sinkc_valid = sinkC_io_resp_valid & _T_18; // @[Scheduler.scala 77:22:chipyard.TestHarness.RocketConfig.fir@100168.4]
  assign abc_mshrs_3_io_sinkc_bits_last = sinkC_io_resp_bits_last; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100175.4]
  assign abc_mshrs_3_io_sinkc_bits_tag = sinkC_io_resp_bits_tag; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100175.4]
  assign abc_mshrs_3_io_sinkc_bits_source = sinkC_io_resp_bits_source; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100175.4]
  assign abc_mshrs_3_io_sinkc_bits_param = sinkC_io_resp_bits_param; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100175.4]
  assign abc_mshrs_3_io_sinkc_bits_data = sinkC_io_resp_bits_data; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100175.4]
  assign abc_mshrs_3_io_sinkd_valid = sinkD_io_resp_valid & _T_20; // @[Scheduler.scala 78:22:chipyard.TestHarness.RocketConfig.fir@100171.4]
  assign abc_mshrs_3_io_sinkd_bits_last = sinkD_io_resp_bits_last; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100176.4]
  assign abc_mshrs_3_io_sinkd_bits_opcode = sinkD_io_resp_bits_opcode; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100176.4]
  assign abc_mshrs_3_io_sinkd_bits_param = sinkD_io_resp_bits_param; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100176.4]
  assign abc_mshrs_3_io_sinkd_bits_sink = sinkD_io_resp_bits_sink; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100176.4]
  assign abc_mshrs_3_io_sinkd_bits_denied = sinkD_io_resp_bits_denied; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100176.4]
  assign abc_mshrs_3_io_sinke_valid = sinkE_io_resp_valid & _T_22; // @[Scheduler.scala 79:22:chipyard.TestHarness.RocketConfig.fir@100174.4]
  assign abc_mshrs_3_io_nestedwb_set = mshr_selectOH[6] ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100178.4]
  assign abc_mshrs_3_io_nestedwb_tag = mshr_selectOH[6] ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100178.4]
  assign abc_mshrs_3_io_nestedwb_b_toN = _T_704 & _T_705; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100178.4]
  assign abc_mshrs_3_io_nestedwb_b_toB = _T_704 & _T_708; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100178.4]
  assign abc_mshrs_3_io_nestedwb_b_clr_dirty = mshr_selectOH[5] & bc_mshr_io_schedule_bits_dir_valid; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100178.4]
  assign abc_mshrs_3_io_nestedwb_c_set_dirty = _T_711 & c_mshr_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100178.4]
  assign abc_mshrs_4_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100115.4]
  assign abc_mshrs_4_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100116.4]
  assign abc_mshrs_4_io_allocate_valid = _T_1194 | _T_987; // @[Scheduler.scala 225:25:chipyard.TestHarness.RocketConfig.fir@101319.4 Scheduler.scala 270:27:chipyard.TestHarness.RocketConfig.fir@101584.6]
  assign abc_mshrs_4_io_allocate_bits_prio_0 = _T_1194 ? request_bits_prio_0 : _T_985_prio_0; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101314.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101585.6]
  assign abc_mshrs_4_io_allocate_bits_prio_1 = _T_1194 ? 1'h0 : _T_985_prio_1; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101314.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101585.6]
  assign abc_mshrs_4_io_allocate_bits_prio_2 = _T_1194 ? request_bits_prio_2 : _T_985_prio_2; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101314.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101585.6]
  assign abc_mshrs_4_io_allocate_bits_control = _T_1194 ? request_bits_control : _T_985_control; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101314.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101585.6]
  assign abc_mshrs_4_io_allocate_bits_opcode = _T_1194 ? request_bits_opcode : _T_985_opcode; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101314.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101585.6]
  assign abc_mshrs_4_io_allocate_bits_param = _T_1194 ? request_bits_param : _T_985_param; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101314.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101585.6]
  assign abc_mshrs_4_io_allocate_bits_size = _T_1194 ? request_bits_size : _T_985_size; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101314.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101585.6]
  assign abc_mshrs_4_io_allocate_bits_source = _T_1194 ? request_bits_source : _T_985_source; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101314.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101585.6]
  assign abc_mshrs_4_io_allocate_bits_tag = _T_1194 ? request_bits_tag : _T_985_tag; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101314.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101585.6]
  assign abc_mshrs_4_io_allocate_bits_offset = _T_1194 ? request_bits_offset : _T_985_offset; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101314.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101585.6]
  assign abc_mshrs_4_io_allocate_bits_put = _T_1194 ? request_bits_put : _T_985_put; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101314.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101585.6]
  assign abc_mshrs_4_io_allocate_bits_set = _T_1194 ? request_bits_set : abc_mshrs_4_io_status_bits_set; // @[Scheduler.scala 223:28:chipyard.TestHarness.RocketConfig.fir@101315.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101585.6]
  assign abc_mshrs_4_io_allocate_bits_repeat = _T_1194 ? 1'h0 : _T_986; // @[Scheduler.scala 224:31:chipyard.TestHarness.RocketConfig.fir@101317.4 Scheduler.scala 272:33:chipyard.TestHarness.RocketConfig.fir@101586.6]
  assign abc_mshrs_4_io_directory_valid = directoryFanout[4]; // @[Scheduler.scala 298:26:chipyard.TestHarness.RocketConfig.fir@101674.4]
  assign abc_mshrs_4_io_directory_bits_dirty = directory_io_result_bits_dirty; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101675.4]
  assign abc_mshrs_4_io_directory_bits_state = directory_io_result_bits_state; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101675.4]
  assign abc_mshrs_4_io_directory_bits_clients = directory_io_result_bits_clients; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101675.4]
  assign abc_mshrs_4_io_directory_bits_tag = directory_io_result_bits_tag; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101675.4]
  assign abc_mshrs_4_io_directory_bits_hit = directory_io_result_bits_hit; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101675.4]
  assign abc_mshrs_4_io_directory_bits_way = directory_io_result_bits_way; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101675.4]
  assign abc_mshrs_4_io_schedule_ready = mshr_selectOH[4]; // @[Scheduler.scala 213:25:chipyard.TestHarness.RocketConfig.fir@101291.4]
  assign abc_mshrs_4_io_sinkc_valid = sinkC_io_resp_valid & _T_24; // @[Scheduler.scala 77:22:chipyard.TestHarness.RocketConfig.fir@100181.4]
  assign abc_mshrs_4_io_sinkc_bits_last = sinkC_io_resp_bits_last; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100188.4]
  assign abc_mshrs_4_io_sinkc_bits_tag = sinkC_io_resp_bits_tag; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100188.4]
  assign abc_mshrs_4_io_sinkc_bits_source = sinkC_io_resp_bits_source; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100188.4]
  assign abc_mshrs_4_io_sinkc_bits_param = sinkC_io_resp_bits_param; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100188.4]
  assign abc_mshrs_4_io_sinkc_bits_data = sinkC_io_resp_bits_data; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100188.4]
  assign abc_mshrs_4_io_sinkd_valid = sinkD_io_resp_valid & _T_26; // @[Scheduler.scala 78:22:chipyard.TestHarness.RocketConfig.fir@100184.4]
  assign abc_mshrs_4_io_sinkd_bits_last = sinkD_io_resp_bits_last; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100189.4]
  assign abc_mshrs_4_io_sinkd_bits_opcode = sinkD_io_resp_bits_opcode; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100189.4]
  assign abc_mshrs_4_io_sinkd_bits_param = sinkD_io_resp_bits_param; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100189.4]
  assign abc_mshrs_4_io_sinkd_bits_sink = sinkD_io_resp_bits_sink; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100189.4]
  assign abc_mshrs_4_io_sinkd_bits_denied = sinkD_io_resp_bits_denied; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100189.4]
  assign abc_mshrs_4_io_sinke_valid = sinkE_io_resp_valid & _T_28; // @[Scheduler.scala 79:22:chipyard.TestHarness.RocketConfig.fir@100187.4]
  assign abc_mshrs_4_io_nestedwb_set = mshr_selectOH[6] ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100191.4]
  assign abc_mshrs_4_io_nestedwb_tag = mshr_selectOH[6] ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100191.4]
  assign abc_mshrs_4_io_nestedwb_b_toN = _T_704 & _T_705; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100191.4]
  assign abc_mshrs_4_io_nestedwb_b_toB = _T_704 & _T_708; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100191.4]
  assign abc_mshrs_4_io_nestedwb_b_clr_dirty = mshr_selectOH[5] & bc_mshr_io_schedule_bits_dir_valid; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100191.4]
  assign abc_mshrs_4_io_nestedwb_c_set_dirty = _T_711 & c_mshr_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100191.4]
  assign bc_mshr_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100119.4]
  assign bc_mshr_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100120.4]
  assign bc_mshr_io_allocate_valid = _T_1198 | _T_1010; // @[Scheduler.scala 225:25:chipyard.TestHarness.RocketConfig.fir@101349.4 Scheduler.scala 270:27:chipyard.TestHarness.RocketConfig.fir@101593.6 Scheduler.scala 277:31:chipyard.TestHarness.RocketConfig.fir@101614.6]
  assign bc_mshr_io_allocate_bits_prio_0 = 1'h0; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101344.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101594.6 Scheduler.scala 278:30:chipyard.TestHarness.RocketConfig.fir@101615.6 Scheduler.scala 282:36:chipyard.TestHarness.RocketConfig.fir@101626.4]
  assign bc_mshr_io_allocate_bits_prio_1 = _T_1198 ? 1'h0 : _T_1008_prio_1; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101344.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101594.6 Scheduler.scala 278:30:chipyard.TestHarness.RocketConfig.fir@101615.6]
  assign bc_mshr_io_allocate_bits_prio_2 = _T_1198 ? request_bits_prio_2 : _T_1008_prio_2; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101344.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101594.6 Scheduler.scala 278:30:chipyard.TestHarness.RocketConfig.fir@101615.6]
  assign bc_mshr_io_allocate_bits_control = _T_1198 ? request_bits_control : _T_1008_control; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101344.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101594.6 Scheduler.scala 278:30:chipyard.TestHarness.RocketConfig.fir@101615.6]
  assign bc_mshr_io_allocate_bits_opcode = _T_1198 ? request_bits_opcode : _T_1008_opcode; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101344.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101594.6 Scheduler.scala 278:30:chipyard.TestHarness.RocketConfig.fir@101615.6]
  assign bc_mshr_io_allocate_bits_param = _T_1198 ? request_bits_param : _T_1008_param; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101344.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101594.6 Scheduler.scala 278:30:chipyard.TestHarness.RocketConfig.fir@101615.6]
  assign bc_mshr_io_allocate_bits_size = _T_1198 ? request_bits_size : _T_1008_size; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101344.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101594.6 Scheduler.scala 278:30:chipyard.TestHarness.RocketConfig.fir@101615.6]
  assign bc_mshr_io_allocate_bits_source = _T_1198 ? request_bits_source : _T_1008_source; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101344.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101594.6 Scheduler.scala 278:30:chipyard.TestHarness.RocketConfig.fir@101615.6]
  assign bc_mshr_io_allocate_bits_tag = _T_1198 ? request_bits_tag : _T_1008_tag; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101344.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101594.6 Scheduler.scala 278:30:chipyard.TestHarness.RocketConfig.fir@101615.6]
  assign bc_mshr_io_allocate_bits_offset = _T_1198 ? request_bits_offset : _T_1008_offset; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101344.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101594.6 Scheduler.scala 278:30:chipyard.TestHarness.RocketConfig.fir@101615.6]
  assign bc_mshr_io_allocate_bits_put = _T_1198 ? request_bits_put : _T_1008_put; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101344.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101594.6 Scheduler.scala 278:30:chipyard.TestHarness.RocketConfig.fir@101615.6]
  assign bc_mshr_io_allocate_bits_set = _T_1198 ? request_bits_set : bc_mshr_io_status_bits_set; // @[Scheduler.scala 223:28:chipyard.TestHarness.RocketConfig.fir@101345.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101594.6 Scheduler.scala 278:30:chipyard.TestHarness.RocketConfig.fir@101615.6]
  assign bc_mshr_io_allocate_bits_repeat = _T_1198 ? 1'h0 : _T_1009; // @[Scheduler.scala 224:31:chipyard.TestHarness.RocketConfig.fir@101347.4 Scheduler.scala 272:33:chipyard.TestHarness.RocketConfig.fir@101595.6 Scheduler.scala 279:37:chipyard.TestHarness.RocketConfig.fir@101616.6]
  assign bc_mshr_io_directory_valid = directoryFanout[5]; // @[Scheduler.scala 298:26:chipyard.TestHarness.RocketConfig.fir@101677.4]
  assign bc_mshr_io_directory_bits_dirty = directory_io_result_bits_dirty; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101678.4]
  assign bc_mshr_io_directory_bits_state = directory_io_result_bits_state; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101678.4]
  assign bc_mshr_io_directory_bits_clients = directory_io_result_bits_clients; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101678.4]
  assign bc_mshr_io_directory_bits_tag = directory_io_result_bits_tag; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101678.4]
  assign bc_mshr_io_directory_bits_hit = directory_io_result_bits_hit; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101678.4]
  assign bc_mshr_io_directory_bits_way = directory_io_result_bits_way; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101678.4]
  assign bc_mshr_io_schedule_ready = mshr_selectOH[5]; // @[Scheduler.scala 213:25:chipyard.TestHarness.RocketConfig.fir@101321.4]
  assign bc_mshr_io_sinkc_valid = sinkC_io_resp_valid & _T_30; // @[Scheduler.scala 77:22:chipyard.TestHarness.RocketConfig.fir@100194.4]
  assign bc_mshr_io_sinkc_bits_last = sinkC_io_resp_bits_last; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100201.4]
  assign bc_mshr_io_sinkc_bits_tag = sinkC_io_resp_bits_tag; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100201.4]
  assign bc_mshr_io_sinkc_bits_source = sinkC_io_resp_bits_source; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100201.4]
  assign bc_mshr_io_sinkc_bits_param = sinkC_io_resp_bits_param; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100201.4]
  assign bc_mshr_io_sinkc_bits_data = sinkC_io_resp_bits_data; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100201.4]
  assign bc_mshr_io_sinkd_valid = sinkD_io_resp_valid & _T_32; // @[Scheduler.scala 78:22:chipyard.TestHarness.RocketConfig.fir@100197.4]
  assign bc_mshr_io_sinkd_bits_last = sinkD_io_resp_bits_last; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100202.4]
  assign bc_mshr_io_sinkd_bits_opcode = sinkD_io_resp_bits_opcode; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100202.4]
  assign bc_mshr_io_sinkd_bits_param = sinkD_io_resp_bits_param; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100202.4]
  assign bc_mshr_io_sinkd_bits_sink = sinkD_io_resp_bits_sink; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100202.4]
  assign bc_mshr_io_sinkd_bits_denied = sinkD_io_resp_bits_denied; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100202.4]
  assign bc_mshr_io_sinke_valid = sinkE_io_resp_valid & _T_34; // @[Scheduler.scala 79:22:chipyard.TestHarness.RocketConfig.fir@100200.4]
  assign bc_mshr_io_nestedwb_set = mshr_selectOH[6] ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100204.4]
  assign bc_mshr_io_nestedwb_tag = mshr_selectOH[6] ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100204.4]
  assign bc_mshr_io_nestedwb_b_toN = _T_704 & _T_705; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100204.4]
  assign bc_mshr_io_nestedwb_b_toB = _T_704 & _T_708; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100204.4]
  assign bc_mshr_io_nestedwb_b_clr_dirty = mshr_selectOH[5] & bc_mshr_io_schedule_bits_dir_valid; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100204.4]
  assign bc_mshr_io_nestedwb_c_set_dirty = _T_711 & c_mshr_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100204.4]
  assign c_mshr_clock = clock; // @[:chipyard.TestHarness.RocketConfig.fir@100123.4]
  assign c_mshr_reset = reset; // @[:chipyard.TestHarness.RocketConfig.fir@100124.4]
  assign c_mshr_io_allocate_valid = _T_1218 | _GEN_85; // @[Scheduler.scala 225:25:chipyard.TestHarness.RocketConfig.fir@101379.4 Scheduler.scala 270:27:chipyard.TestHarness.RocketConfig.fir@101602.6 Scheduler.scala 285:30:chipyard.TestHarness.RocketConfig.fir@101633.6]
  assign c_mshr_io_allocate_bits_prio_0 = 1'h0; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101374.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101603.6 Scheduler.scala 286:29:chipyard.TestHarness.RocketConfig.fir@101634.6 Scheduler.scala 291:35:chipyard.TestHarness.RocketConfig.fir@101653.4]
  assign c_mshr_io_allocate_bits_prio_1 = 1'h0; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101374.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101603.6 Scheduler.scala 286:29:chipyard.TestHarness.RocketConfig.fir@101634.6 Scheduler.scala 292:35:chipyard.TestHarness.RocketConfig.fir@101654.4]
  assign c_mshr_io_allocate_bits_prio_2 = _T_1218 ? request_bits_prio_2 : _GEN_88; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101374.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101603.6 Scheduler.scala 286:29:chipyard.TestHarness.RocketConfig.fir@101634.6]
  assign c_mshr_io_allocate_bits_control = _T_1218 ? request_bits_control : _GEN_89; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101374.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101603.6 Scheduler.scala 286:29:chipyard.TestHarness.RocketConfig.fir@101634.6]
  assign c_mshr_io_allocate_bits_opcode = _T_1218 ? request_bits_opcode : _GEN_90; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101374.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101603.6 Scheduler.scala 286:29:chipyard.TestHarness.RocketConfig.fir@101634.6]
  assign c_mshr_io_allocate_bits_param = _T_1218 ? request_bits_param : _GEN_91; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101374.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101603.6 Scheduler.scala 286:29:chipyard.TestHarness.RocketConfig.fir@101634.6]
  assign c_mshr_io_allocate_bits_size = _T_1218 ? request_bits_size : _GEN_92; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101374.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101603.6 Scheduler.scala 286:29:chipyard.TestHarness.RocketConfig.fir@101634.6]
  assign c_mshr_io_allocate_bits_source = _T_1218 ? request_bits_source : _GEN_93; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101374.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101603.6 Scheduler.scala 286:29:chipyard.TestHarness.RocketConfig.fir@101634.6]
  assign c_mshr_io_allocate_bits_tag = _T_1218 ? request_bits_tag : _GEN_94; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101374.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101603.6 Scheduler.scala 286:29:chipyard.TestHarness.RocketConfig.fir@101634.6]
  assign c_mshr_io_allocate_bits_offset = _T_1218 ? request_bits_offset : _GEN_95; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101374.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101603.6 Scheduler.scala 286:29:chipyard.TestHarness.RocketConfig.fir@101634.6]
  assign c_mshr_io_allocate_bits_put = _T_1218 ? request_bits_put : _GEN_96; // @[Scheduler.scala 222:24:chipyard.TestHarness.RocketConfig.fir@101374.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101603.6 Scheduler.scala 286:29:chipyard.TestHarness.RocketConfig.fir@101634.6]
  assign c_mshr_io_allocate_bits_set = _T_1218 ? request_bits_set : _GEN_97; // @[Scheduler.scala 223:28:chipyard.TestHarness.RocketConfig.fir@101375.4 Scheduler.scala 271:26:chipyard.TestHarness.RocketConfig.fir@101603.6 Scheduler.scala 286:29:chipyard.TestHarness.RocketConfig.fir@101634.6]
  assign c_mshr_io_allocate_bits_repeat = _T_1218 ? 1'h0 : _GEN_98; // @[Scheduler.scala 224:31:chipyard.TestHarness.RocketConfig.fir@101377.4 Scheduler.scala 272:33:chipyard.TestHarness.RocketConfig.fir@101604.6 Scheduler.scala 287:36:chipyard.TestHarness.RocketConfig.fir@101635.6]
  assign c_mshr_io_directory_valid = directoryFanout[6]; // @[Scheduler.scala 298:26:chipyard.TestHarness.RocketConfig.fir@101680.4]
  assign c_mshr_io_directory_bits_dirty = directory_io_result_bits_dirty; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101681.4]
  assign c_mshr_io_directory_bits_state = directory_io_result_bits_state; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101681.4]
  assign c_mshr_io_directory_bits_clients = directory_io_result_bits_clients; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101681.4]
  assign c_mshr_io_directory_bits_tag = directory_io_result_bits_tag; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101681.4]
  assign c_mshr_io_directory_bits_hit = directory_io_result_bits_hit; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101681.4]
  assign c_mshr_io_directory_bits_way = directory_io_result_bits_way; // @[Scheduler.scala 299:25:chipyard.TestHarness.RocketConfig.fir@101681.4]
  assign c_mshr_io_schedule_ready = mshr_selectOH[6]; // @[Scheduler.scala 213:25:chipyard.TestHarness.RocketConfig.fir@101351.4]
  assign c_mshr_io_sinkc_valid = sinkC_io_resp_valid & _T_36; // @[Scheduler.scala 77:22:chipyard.TestHarness.RocketConfig.fir@100207.4]
  assign c_mshr_io_sinkc_bits_last = sinkC_io_resp_bits_last; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100214.4]
  assign c_mshr_io_sinkc_bits_tag = sinkC_io_resp_bits_tag; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100214.4]
  assign c_mshr_io_sinkc_bits_source = sinkC_io_resp_bits_source; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100214.4]
  assign c_mshr_io_sinkc_bits_param = sinkC_io_resp_bits_param; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100214.4]
  assign c_mshr_io_sinkc_bits_data = sinkC_io_resp_bits_data; // @[Scheduler.scala 80:21:chipyard.TestHarness.RocketConfig.fir@100214.4]
  assign c_mshr_io_sinkd_valid = sinkD_io_resp_valid & _T_38; // @[Scheduler.scala 78:22:chipyard.TestHarness.RocketConfig.fir@100210.4]
  assign c_mshr_io_sinkd_bits_last = sinkD_io_resp_bits_last; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100215.4]
  assign c_mshr_io_sinkd_bits_opcode = sinkD_io_resp_bits_opcode; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100215.4]
  assign c_mshr_io_sinkd_bits_param = sinkD_io_resp_bits_param; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100215.4]
  assign c_mshr_io_sinkd_bits_sink = sinkD_io_resp_bits_sink; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100215.4]
  assign c_mshr_io_sinkd_bits_denied = sinkD_io_resp_bits_denied; // @[Scheduler.scala 81:21:chipyard.TestHarness.RocketConfig.fir@100215.4]
  assign c_mshr_io_sinke_valid = sinkE_io_resp_valid & _T_40; // @[Scheduler.scala 79:22:chipyard.TestHarness.RocketConfig.fir@100213.4]
  assign c_mshr_io_nestedwb_set = mshr_selectOH[6] ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100217.4]
  assign c_mshr_io_nestedwb_tag = mshr_selectOH[6] ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100217.4]
  assign c_mshr_io_nestedwb_b_toN = _T_704 & _T_705; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100217.4]
  assign c_mshr_io_nestedwb_b_toB = _T_704 & _T_708; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100217.4]
  assign c_mshr_io_nestedwb_b_clr_dirty = mshr_selectOH[5] & bc_mshr_io_schedule_bits_dir_valid; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100217.4]
  assign c_mshr_io_nestedwb_c_set_dirty = _T_711 & c_mshr_io_schedule_bits_dir_bits_data_dirty; // @[Scheduler.scala 83:19:chipyard.TestHarness.RocketConfig.fir@100217.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  robin_filter = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  directoryFanout = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      robin_filter <= 7'h0;
    end else if (_T_691) begin
      robin_filter <= _T_699;
    end
    if (mshr_uses_directory) begin
      directoryFanout <= {{1'd0}, mshr_selectOH};
    end else if (alloc_uses_directory) begin
      if (alloc) begin
        directoryFanout <= mshr_insertOH;
      end else begin
        directoryFanout <= 8'h40;
      end
    end else begin
      directoryFanout <= 8'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1218 & _T_1213) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Scheduler.scala:288 assert (!request.bits.prio(0))\n"); // @[Scheduler.scala 288:12:chipyard.TestHarness.RocketConfig.fir@101641.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1218 & _T_1213) begin
          $fatal; // @[Scheduler.scala 288:12:chipyard.TestHarness.RocketConfig.fir@101642.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
