module FPUDecoder( // @[:chipyard.TestHarness.RocketConfig.fir@233345.2]
  input  [31:0] io_inst, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_wen, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_ren1, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_ren2, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_ren3, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_swap12, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_swap23, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_singleIn, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_singleOut, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_fromint, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_toint, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_fastpipe, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_fma, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_div, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_sqrt, // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
  output        io_sigs_wflags // @[:chipyard.TestHarness.RocketConfig.fir@233348.4]
);
  wire [31:0] _T; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233353.4]
  wire [31:0] _T_2; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233356.4]
  wire  _T_3; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233357.4]
  wire [31:0] _T_4; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233358.4]
  wire  _T_5; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233359.4]
  wire [31:0] _T_6; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233360.4]
  wire  _T_7; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233361.4]
  wire  _T_9; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233363.4]
  wire [31:0] _T_10; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233365.4]
  wire  _T_11; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233366.4]
  wire [31:0] _T_12; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233367.4]
  wire  _T_13; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233368.4]
  wire [31:0] _T_14; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233369.4]
  wire  decoder_4; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233370.4]
  wire  _T_17; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233372.4]
  wire [31:0] _T_18; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233374.4]
  wire  _T_19; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233375.4]
  wire [31:0] _T_20; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233376.4]
  wire  _T_21; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233377.4]
  wire  _T_23; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233379.4]
  wire [31:0] _T_24; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233383.4]
  wire [31:0] _T_26; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233386.4]
  wire  _T_27; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233387.4]
  wire [31:0] _T_28; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233388.4]
  wire  _T_29; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233389.4]
  wire [31:0] _T_30; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233390.4]
  wire  _T_31; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233391.4]
  wire [31:0] _T_32; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233392.4]
  wire  _T_33; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233393.4]
  wire [31:0] _T_34; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233394.4]
  wire  _T_35; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233395.4]
  wire [31:0] _T_36; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233396.4]
  wire  _T_37; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233397.4]
  wire [31:0] _T_38; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233398.4]
  wire  _T_39; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233399.4]
  wire  _T_41; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233401.4]
  wire  _T_42; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233402.4]
  wire  _T_43; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233403.4]
  wire  _T_44; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233404.4]
  wire  _T_45; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233405.4]
  wire [31:0] _T_46; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233407.4]
  wire  _T_47; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233408.4]
  wire [31:0] _T_48; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233409.4]
  wire  _T_49; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233410.4]
  wire  _T_51; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233412.4]
  wire [31:0] _T_52; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233413.4]
  wire  _T_53; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233414.4]
  wire [31:0] _T_54; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233415.4]
  wire  _T_55; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233416.4]
  wire  _T_57; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233418.4]
  wire  _T_58; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233419.4]
  wire  _T_59; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233420.4]
  wire [31:0] _T_60; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233422.4]
  wire  _T_63; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233426.4]
  wire [31:0] _T_65; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233429.4]
  wire  _T_66; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233430.4]
  wire [31:0] _T_67; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233431.4]
  wire  _T_68; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233432.4]
  wire [31:0] _T_70; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233435.4]
  wire  _T_71; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233436.4]
  wire [31:0] _T_72; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233437.4]
  wire  _T_73; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233438.4]
  wire  _T_75; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233440.4]
  wire [31:0] _T_76; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233442.4]
  wire [31:0] _T_80; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233448.4]
  wire  _T_81; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233449.4]
  wire [31:0] _T_82; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233450.4]
  wire  _T_83; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233451.4]
  wire [31:0] _T_84; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233452.4]
  wire  _T_85; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233453.4]
  wire  _T_87; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233455.4]
  wire  _T_88; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233456.4]
  assign _T = io_inst & 32'h40; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233353.4]
  assign _T_2 = io_inst & 32'h80000020; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233356.4]
  assign _T_3 = _T_2 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233357.4]
  assign _T_4 = io_inst & 32'h30; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233358.4]
  assign _T_5 = _T_4 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233359.4]
  assign _T_6 = io_inst & 32'h10000020; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233360.4]
  assign _T_7 = _T_6 == 32'h10000000; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233361.4]
  assign _T_9 = _T_3 | _T_5; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233363.4]
  assign _T_10 = io_inst & 32'h80000004; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233365.4]
  assign _T_11 = _T_10 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233366.4]
  assign _T_12 = io_inst & 32'h10000004; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233367.4]
  assign _T_13 = _T_12 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233368.4]
  assign _T_14 = io_inst & 32'h50; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233369.4]
  assign decoder_4 = _T_14 == 32'h40; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233370.4]
  assign _T_17 = _T_11 | _T_13; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233372.4]
  assign _T_18 = io_inst & 32'h40000004; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233374.4]
  assign _T_19 = _T_18 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233375.4]
  assign _T_20 = io_inst & 32'h20; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233376.4]
  assign _T_21 = _T_20 == 32'h20; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233377.4]
  assign _T_23 = _T_19 | _T_21; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233379.4]
  assign _T_24 = io_inst & 32'h30000010; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233383.4]
  assign _T_26 = io_inst & 32'h82100020; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233386.4]
  assign _T_27 = _T_26 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233387.4]
  assign _T_28 = io_inst & 32'h42000020; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233388.4]
  assign _T_29 = _T_28 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233389.4]
  assign _T_30 = io_inst & 32'h2000030; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233390.4]
  assign _T_31 = _T_30 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233391.4]
  assign _T_32 = io_inst & 32'h2103000; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233392.4]
  assign _T_33 = _T_32 == 32'h1000; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233393.4]
  assign _T_34 = io_inst & 32'h12002000; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233394.4]
  assign _T_35 = _T_34 == 32'h10000000; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233395.4]
  assign _T_36 = io_inst & 32'hd0100010; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233396.4]
  assign _T_37 = _T_36 == 32'h40000010; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233397.4]
  assign _T_38 = io_inst & 32'ha2000020; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233398.4]
  assign _T_39 = _T_38 == 32'h80000000; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233399.4]
  assign _T_41 = _T_27 | _T_29; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233401.4]
  assign _T_42 = _T_41 | _T_31; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233402.4]
  assign _T_43 = _T_42 | _T_33; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233403.4]
  assign _T_44 = _T_43 | _T_35; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233404.4]
  assign _T_45 = _T_44 | _T_37; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233405.4]
  assign _T_46 = io_inst & 32'h42001000; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233407.4]
  assign _T_47 = _T_46 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233408.4]
  assign _T_48 = io_inst & 32'h22000004; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233409.4]
  assign _T_49 = _T_48 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233410.4]
  assign _T_51 = _T_34 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233412.4]
  assign _T_52 = io_inst & 32'h1040; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233413.4]
  assign _T_53 = _T_52 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233414.4]
  assign _T_54 = io_inst & 32'h2000050; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233415.4]
  assign _T_55 = _T_54 == 32'h40; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233416.4]
  assign _T_57 = _T_47 | _T_49; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233418.4]
  assign _T_58 = _T_57 | _T_51; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233419.4]
  assign _T_59 = _T_58 | _T_53; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233420.4]
  assign _T_60 = io_inst & 32'h90000010; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233422.4]
  assign _T_63 = _T_60 == 32'h80000010; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233426.4]
  assign _T_65 = io_inst & 32'ha0000010; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233429.4]
  assign _T_66 = _T_65 == 32'h20000010; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233430.4]
  assign _T_67 = io_inst & 32'hd0000010; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233431.4]
  assign _T_68 = _T_67 == 32'h40000010; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233432.4]
  assign _T_70 = io_inst & 32'h70000004; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233435.4]
  assign _T_71 = _T_70 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233436.4]
  assign _T_72 = io_inst & 32'h68000004; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233437.4]
  assign _T_73 = _T_72 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233438.4]
  assign _T_75 = _T_71 | _T_73; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233440.4]
  assign _T_76 = io_inst & 32'h58000010; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233442.4]
  assign _T_80 = io_inst & 32'h20000004; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233448.4]
  assign _T_81 = _T_80 == 32'h0; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233449.4]
  assign _T_82 = io_inst & 32'h8002000; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233450.4]
  assign _T_83 = _T_82 == 32'h8000000; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233451.4]
  assign _T_84 = io_inst & 32'hc0000004; // @[Decode.scala 14:65:chipyard.TestHarness.RocketConfig.fir@233452.4]
  assign _T_85 = _T_84 == 32'h80000000; // @[Decode.scala 14:121:chipyard.TestHarness.RocketConfig.fir@233453.4]
  assign _T_87 = _T_81 | decoder_4; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233455.4]
  assign _T_88 = _T_87 | _T_83; // @[Decode.scala 15:30:chipyard.TestHarness.RocketConfig.fir@233456.4]
  assign io_sigs_wen = _T_9 | _T_7; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233459.4]
  assign io_sigs_ren1 = _T_17 | decoder_4; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233460.4]
  assign io_sigs_ren2 = _T_23 | decoder_4; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233461.4]
  assign io_sigs_ren3 = _T_14 == 32'h40; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233462.4]
  assign io_sigs_swap12 = _T == 32'h0; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233463.4]
  assign io_sigs_swap23 = _T_24 == 32'h10; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233464.4]
  assign io_sigs_singleIn = _T_45 | _T_39; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233465.4]
  assign io_sigs_singleOut = _T_59 | _T_55; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233466.4]
  assign io_sigs_fromint = _T_60 == 32'h90000010; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233467.4]
  assign io_sigs_toint = _T_21 | _T_63; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233468.4]
  assign io_sigs_fastpipe = _T_66 | _T_68; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233469.4]
  assign io_sigs_fma = _T_75 | decoder_4; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233470.4]
  assign io_sigs_div = _T_76 == 32'h18000010; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233471.4]
  assign io_sigs_sqrt = _T_67 == 32'h50000010; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233472.4]
  assign io_sigs_wflags = _T_88 | _T_85; // @[FPU.scala 135:40:chipyard.TestHarness.RocketConfig.fir@233473.4]
endmodule
