module MSHR( // @[:chipyard.TestHarness.RocketConfig.fir@89164.2]
  input         clock, // @[:chipyard.TestHarness.RocketConfig.fir@89165.4]
  input         reset, // @[:chipyard.TestHarness.RocketConfig.fir@89166.4]
  input         io_allocate_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_allocate_bits_prio_0, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_allocate_bits_prio_1, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_allocate_bits_prio_2, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_allocate_bits_control, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [2:0]  io_allocate_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [2:0]  io_allocate_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [2:0]  io_allocate_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [2:0]  io_allocate_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [11:0] io_allocate_bits_tag, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [5:0]  io_allocate_bits_offset, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [5:0]  io_allocate_bits_put, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [9:0]  io_allocate_bits_set, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_allocate_bits_repeat, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_directory_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_directory_bits_dirty, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [1:0]  io_directory_bits_state, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_directory_bits_clients, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [11:0] io_directory_bits_tag, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_directory_bits_hit, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [2:0]  io_directory_bits_way, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_status_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [9:0]  io_status_bits_set, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [11:0] io_status_bits_tag, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [2:0]  io_status_bits_way, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_status_bits_blockB, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_status_bits_nestB, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_status_bits_blockC, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_status_bits_nestC, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_schedule_ready, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_a_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [11:0] io_schedule_bits_a_bits_tag, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [9:0]  io_schedule_bits_a_bits_set, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [2:0]  io_schedule_bits_a_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_a_bits_block, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_b_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [2:0]  io_schedule_bits_b_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [11:0] io_schedule_bits_b_bits_tag, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [9:0]  io_schedule_bits_b_bits_set, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_b_bits_clients, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_c_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [2:0]  io_schedule_bits_c_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [2:0]  io_schedule_bits_c_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [11:0] io_schedule_bits_c_bits_tag, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [9:0]  io_schedule_bits_c_bits_set, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [2:0]  io_schedule_bits_c_bits_way, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_c_bits_dirty, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_d_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_d_bits_prio_0, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_d_bits_prio_1, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_d_bits_prio_2, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_d_bits_control, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [2:0]  io_schedule_bits_d_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [2:0]  io_schedule_bits_d_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [2:0]  io_schedule_bits_d_bits_size, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [2:0]  io_schedule_bits_d_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [11:0] io_schedule_bits_d_bits_tag, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [5:0]  io_schedule_bits_d_bits_offset, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [5:0]  io_schedule_bits_d_bits_put, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [9:0]  io_schedule_bits_d_bits_set, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [2:0]  io_schedule_bits_d_bits_way, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_d_bits_bad, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_e_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [2:0]  io_schedule_bits_e_bits_sink, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_x_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_dir_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [9:0]  io_schedule_bits_dir_bits_set, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [2:0]  io_schedule_bits_dir_bits_way, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_dir_bits_data_dirty, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [1:0]  io_schedule_bits_dir_bits_data_state, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_dir_bits_data_clients, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output [11:0] io_schedule_bits_dir_bits_data_tag, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  output        io_schedule_bits_reload, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_sinkc_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_sinkc_bits_last, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [11:0] io_sinkc_bits_tag, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [2:0]  io_sinkc_bits_source, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [2:0]  io_sinkc_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_sinkc_bits_data, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_sinkd_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_sinkd_bits_last, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [2:0]  io_sinkd_bits_opcode, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [2:0]  io_sinkd_bits_param, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [2:0]  io_sinkd_bits_sink, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_sinkd_bits_denied, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_sinke_valid, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [9:0]  io_nestedwb_set, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input  [11:0] io_nestedwb_tag, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_nestedwb_b_toN, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_nestedwb_b_toB, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_nestedwb_b_clr_dirty, // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
  input         io_nestedwb_c_set_dirty // @[:chipyard.TestHarness.RocketConfig.fir@89167.4]
);
  reg  request_valid; // @[MSHR.scala 94:30:chipyard.TestHarness.RocketConfig.fir@89172.4]
  reg [31:0] _RAND_0;
  reg  request_prio_0; // @[MSHR.scala 95:20:chipyard.TestHarness.RocketConfig.fir@89173.4]
  reg [31:0] _RAND_1;
  reg  request_prio_1; // @[MSHR.scala 95:20:chipyard.TestHarness.RocketConfig.fir@89173.4]
  reg [31:0] _RAND_2;
  reg  request_prio_2; // @[MSHR.scala 95:20:chipyard.TestHarness.RocketConfig.fir@89173.4]
  reg [31:0] _RAND_3;
  reg  request_control; // @[MSHR.scala 95:20:chipyard.TestHarness.RocketConfig.fir@89173.4]
  reg [31:0] _RAND_4;
  reg [2:0] request_opcode; // @[MSHR.scala 95:20:chipyard.TestHarness.RocketConfig.fir@89173.4]
  reg [31:0] _RAND_5;
  reg [2:0] request_param; // @[MSHR.scala 95:20:chipyard.TestHarness.RocketConfig.fir@89173.4]
  reg [31:0] _RAND_6;
  reg [2:0] request_size; // @[MSHR.scala 95:20:chipyard.TestHarness.RocketConfig.fir@89173.4]
  reg [31:0] _RAND_7;
  reg [2:0] request_source; // @[MSHR.scala 95:20:chipyard.TestHarness.RocketConfig.fir@89173.4]
  reg [31:0] _RAND_8;
  reg [11:0] request_tag; // @[MSHR.scala 95:20:chipyard.TestHarness.RocketConfig.fir@89173.4]
  reg [31:0] _RAND_9;
  reg [5:0] request_offset; // @[MSHR.scala 95:20:chipyard.TestHarness.RocketConfig.fir@89173.4]
  reg [31:0] _RAND_10;
  reg [5:0] request_put; // @[MSHR.scala 95:20:chipyard.TestHarness.RocketConfig.fir@89173.4]
  reg [31:0] _RAND_11;
  reg [9:0] request_set; // @[MSHR.scala 95:20:chipyard.TestHarness.RocketConfig.fir@89173.4]
  reg [31:0] _RAND_12;
  reg  meta_valid; // @[MSHR.scala 96:27:chipyard.TestHarness.RocketConfig.fir@89174.4]
  reg [31:0] _RAND_13;
  reg  meta_dirty; // @[MSHR.scala 97:17:chipyard.TestHarness.RocketConfig.fir@89175.4]
  reg [31:0] _RAND_14;
  reg [1:0] meta_state; // @[MSHR.scala 97:17:chipyard.TestHarness.RocketConfig.fir@89175.4]
  reg [31:0] _RAND_15;
  reg  meta_clients; // @[MSHR.scala 97:17:chipyard.TestHarness.RocketConfig.fir@89175.4]
  reg [31:0] _RAND_16;
  reg [11:0] meta_tag; // @[MSHR.scala 97:17:chipyard.TestHarness.RocketConfig.fir@89175.4]
  reg [31:0] _RAND_17;
  reg  meta_hit; // @[MSHR.scala 97:17:chipyard.TestHarness.RocketConfig.fir@89175.4]
  reg [31:0] _RAND_18;
  reg [2:0] meta_way; // @[MSHR.scala 97:17:chipyard.TestHarness.RocketConfig.fir@89175.4]
  reg [31:0] _RAND_19;
  wire  _T; // @[MSHR.scala 101:22:chipyard.TestHarness.RocketConfig.fir@89177.6]
  wire  _T_1; // @[MSHR.scala 102:29:chipyard.TestHarness.RocketConfig.fir@89179.8]
  wire  _T_2; // @[MSHR.scala 102:15:chipyard.TestHarness.RocketConfig.fir@89180.8]
  wire  _T_4; // @[MSHR.scala 102:14:chipyard.TestHarness.RocketConfig.fir@89182.8]
  wire  _T_5; // @[MSHR.scala 102:14:chipyard.TestHarness.RocketConfig.fir@89183.8]
  wire  _T_6; // @[MSHR.scala 103:15:chipyard.TestHarness.RocketConfig.fir@89188.8]
  wire  _T_8; // @[MSHR.scala 103:14:chipyard.TestHarness.RocketConfig.fir@89190.8]
  wire  _T_9; // @[MSHR.scala 103:14:chipyard.TestHarness.RocketConfig.fir@89191.8]
  wire  _T_10; // @[MSHR.scala 105:22:chipyard.TestHarness.RocketConfig.fir@89197.6]
  wire  _T_15; // @[MSHR.scala 108:22:chipyard.TestHarness.RocketConfig.fir@89208.6]
  wire  _T_18; // @[MSHR.scala 109:14:chipyard.TestHarness.RocketConfig.fir@89212.8]
  wire  _T_19; // @[MSHR.scala 109:14:chipyard.TestHarness.RocketConfig.fir@89213.8]
  wire  _T_21; // @[MSHR.scala 110:45:chipyard.TestHarness.RocketConfig.fir@89219.8]
  wire  _T_22; // @[MSHR.scala 110:29:chipyard.TestHarness.RocketConfig.fir@89220.8]
  wire  _T_23; // @[MSHR.scala 110:57:chipyard.TestHarness.RocketConfig.fir@89221.8]
  wire  _T_25; // @[MSHR.scala 110:14:chipyard.TestHarness.RocketConfig.fir@89223.8]
  wire  _T_26; // @[MSHR.scala 110:14:chipyard.TestHarness.RocketConfig.fir@89224.8]
  wire  _T_27; // @[MSHR.scala 112:22:chipyard.TestHarness.RocketConfig.fir@89230.6]
  reg  s_rprobe; // @[MSHR.scala 118:33:chipyard.TestHarness.RocketConfig.fir@89234.4]
  reg [31:0] _RAND_20;
  reg  w_rprobeackfirst; // @[MSHR.scala 119:33:chipyard.TestHarness.RocketConfig.fir@89235.4]
  reg [31:0] _RAND_21;
  reg  w_rprobeacklast; // @[MSHR.scala 120:33:chipyard.TestHarness.RocketConfig.fir@89236.4]
  reg [31:0] _RAND_22;
  reg  s_release; // @[MSHR.scala 121:33:chipyard.TestHarness.RocketConfig.fir@89237.4]
  reg [31:0] _RAND_23;
  reg  w_releaseack; // @[MSHR.scala 122:33:chipyard.TestHarness.RocketConfig.fir@89238.4]
  reg [31:0] _RAND_24;
  reg  s_pprobe; // @[MSHR.scala 123:33:chipyard.TestHarness.RocketConfig.fir@89239.4]
  reg [31:0] _RAND_25;
  reg  s_acquire; // @[MSHR.scala 124:33:chipyard.TestHarness.RocketConfig.fir@89240.4]
  reg [31:0] _RAND_26;
  reg  s_flush; // @[MSHR.scala 125:33:chipyard.TestHarness.RocketConfig.fir@89241.4]
  reg [31:0] _RAND_27;
  reg  w_grantfirst; // @[MSHR.scala 126:33:chipyard.TestHarness.RocketConfig.fir@89242.4]
  reg [31:0] _RAND_28;
  reg  w_grantlast; // @[MSHR.scala 127:33:chipyard.TestHarness.RocketConfig.fir@89243.4]
  reg [31:0] _RAND_29;
  reg  w_grant; // @[MSHR.scala 128:33:chipyard.TestHarness.RocketConfig.fir@89244.4]
  reg [31:0] _RAND_30;
  reg  w_pprobeackfirst; // @[MSHR.scala 129:33:chipyard.TestHarness.RocketConfig.fir@89245.4]
  reg [31:0] _RAND_31;
  reg  w_pprobeacklast; // @[MSHR.scala 130:33:chipyard.TestHarness.RocketConfig.fir@89246.4]
  reg [31:0] _RAND_32;
  reg  w_pprobeack; // @[MSHR.scala 131:33:chipyard.TestHarness.RocketConfig.fir@89247.4]
  reg [31:0] _RAND_33;
  reg  s_grantack; // @[MSHR.scala 133:33:chipyard.TestHarness.RocketConfig.fir@89249.4]
  reg [31:0] _RAND_34;
  reg  s_execute; // @[MSHR.scala 134:33:chipyard.TestHarness.RocketConfig.fir@89250.4]
  reg [31:0] _RAND_35;
  reg  w_grantack; // @[MSHR.scala 135:33:chipyard.TestHarness.RocketConfig.fir@89251.4]
  reg [31:0] _RAND_36;
  reg  s_writeback; // @[MSHR.scala 136:33:chipyard.TestHarness.RocketConfig.fir@89252.4]
  reg [31:0] _RAND_37;
  reg [2:0] sink; // @[MSHR.scala 144:17:chipyard.TestHarness.RocketConfig.fir@89253.4]
  reg [31:0] _RAND_38;
  reg  gotT; // @[MSHR.scala 145:17:chipyard.TestHarness.RocketConfig.fir@89254.4]
  reg [31:0] _RAND_39;
  reg  bad_grant; // @[MSHR.scala 146:22:chipyard.TestHarness.RocketConfig.fir@89255.4]
  reg [31:0] _RAND_40;
  reg  probes_done; // @[MSHR.scala 147:24:chipyard.TestHarness.RocketConfig.fir@89256.4]
  reg [31:0] _RAND_41;
  reg  probes_toN; // @[MSHR.scala 148:23:chipyard.TestHarness.RocketConfig.fir@89257.4]
  reg [31:0] _RAND_42;
  wire  _T_28; // @[MSHR.scala 152:34:chipyard.TestHarness.RocketConfig.fir@89259.4]
  wire  _T_29; // @[MSHR.scala 152:20:chipyard.TestHarness.RocketConfig.fir@89260.4]
  wire  _T_30; // @[MSHR.scala 153:25:chipyard.TestHarness.RocketConfig.fir@89261.4]
  wire  _T_31; // @[MSHR.scala 152:46:chipyard.TestHarness.RocketConfig.fir@89262.4]
  wire  _T_32; // @[MSHR.scala 153:60:chipyard.TestHarness.RocketConfig.fir@89263.4]
  wire  _T_33; // @[MSHR.scala 153:41:chipyard.TestHarness.RocketConfig.fir@89264.4]
  wire  _GEN_0; // @[MSHR.scala 154:36:chipyard.TestHarness.RocketConfig.fir@89266.6]
  wire  _GEN_1; // @[MSHR.scala 155:36:chipyard.TestHarness.RocketConfig.fir@89269.6]
  wire  _GEN_4; // @[MSHR.scala 153:74:chipyard.TestHarness.RocketConfig.fir@89265.4]
  wire  _T_34; // @[MSHR.scala 165:28:chipyard.TestHarness.RocketConfig.fir@89283.4]
  wire  _T_35; // @[MSHR.scala 165:45:chipyard.TestHarness.RocketConfig.fir@89284.4]
  wire  _T_36; // @[MSHR.scala 165:62:chipyard.TestHarness.RocketConfig.fir@89285.4]
  wire  _T_37; // @[MSHR.scala 165:59:chipyard.TestHarness.RocketConfig.fir@89286.4]
  wire  _T_38; // @[MSHR.scala 165:82:chipyard.TestHarness.RocketConfig.fir@89287.4]
  wire  _T_39; // @[MSHR.scala 165:79:chipyard.TestHarness.RocketConfig.fir@89288.4]
  wire  _T_40; // @[MSHR.scala 165:103:chipyard.TestHarness.RocketConfig.fir@89289.4]
  wire  _T_41; // @[MSHR.scala 165:100:chipyard.TestHarness.RocketConfig.fir@89290.4]
  wire  _T_43; // @[MSHR.scala 166:39:chipyard.TestHarness.RocketConfig.fir@89293.4]
  wire  _T_44; // @[MSHR.scala 166:55:chipyard.TestHarness.RocketConfig.fir@89294.4]
  wire  _T_45; // @[MSHR.scala 166:74:chipyard.TestHarness.RocketConfig.fir@89295.4]
  wire  _T_49; // @[MSHR.scala 170:43:chipyard.TestHarness.RocketConfig.fir@89301.4]
  wire  _T_50; // @[MSHR.scala 170:64:chipyard.TestHarness.RocketConfig.fir@89302.4]
  wire  _T_51; // @[MSHR.scala 170:61:chipyard.TestHarness.RocketConfig.fir@89303.4]
  wire  _T_53; // @[MSHR.scala 170:82:chipyard.TestHarness.RocketConfig.fir@89305.4]
  wire  _T_55; // @[MSHR.scala 176:11:chipyard.TestHarness.RocketConfig.fir@89308.4]
  wire  _T_56; // @[MSHR.scala 176:36:chipyard.TestHarness.RocketConfig.fir@89309.4]
  wire  _T_57; // @[MSHR.scala 176:33:chipyard.TestHarness.RocketConfig.fir@89310.4]
  wire  _T_59; // @[MSHR.scala 176:10:chipyard.TestHarness.RocketConfig.fir@89312.4]
  wire  _T_60; // @[MSHR.scala 176:10:chipyard.TestHarness.RocketConfig.fir@89313.4]
  wire  _T_61; // @[MSHR.scala 177:11:chipyard.TestHarness.RocketConfig.fir@89318.4]
  wire  _T_62; // @[MSHR.scala 177:36:chipyard.TestHarness.RocketConfig.fir@89319.4]
  wire  _T_63; // @[MSHR.scala 177:33:chipyard.TestHarness.RocketConfig.fir@89320.4]
  wire  _T_65; // @[MSHR.scala 177:10:chipyard.TestHarness.RocketConfig.fir@89322.4]
  wire  _T_66; // @[MSHR.scala 177:10:chipyard.TestHarness.RocketConfig.fir@89323.4]
  wire  _T_67; // @[MSHR.scala 180:33:chipyard.TestHarness.RocketConfig.fir@89328.4]
  wire  _T_68; // @[MSHR.scala 180:49:chipyard.TestHarness.RocketConfig.fir@89329.4]
  wire  _T_69; // @[MSHR.scala 180:64:chipyard.TestHarness.RocketConfig.fir@89330.4]
  wire  no_wait; // @[MSHR.scala 180:83:chipyard.TestHarness.RocketConfig.fir@89331.4]
  wire  _T_70; // @[MSHR.scala 181:31:chipyard.TestHarness.RocketConfig.fir@89332.4]
  wire  _T_71; // @[MSHR.scala 181:42:chipyard.TestHarness.RocketConfig.fir@89333.4]
  wire  _T_73; // @[MSHR.scala 182:31:chipyard.TestHarness.RocketConfig.fir@89336.4]
  wire  _T_74; // @[MSHR.scala 182:44:chipyard.TestHarness.RocketConfig.fir@89337.4]
  wire  _T_76; // @[MSHR.scala 183:32:chipyard.TestHarness.RocketConfig.fir@89340.4]
  wire  _T_77; // @[MSHR.scala 183:43:chipyard.TestHarness.RocketConfig.fir@89341.4]
  wire  _T_81; // @[MSHR.scala 184:31:chipyard.TestHarness.RocketConfig.fir@89346.4]
  wire  _T_82; // @[MSHR.scala 184:42:chipyard.TestHarness.RocketConfig.fir@89347.4]
  wire  _T_84; // @[MSHR.scala 185:31:chipyard.TestHarness.RocketConfig.fir@89350.4]
  wire  _T_86; // @[MSHR.scala 186:31:chipyard.TestHarness.RocketConfig.fir@89353.4]
  wire  _T_90; // @[MSHR.scala 187:70:chipyard.TestHarness.RocketConfig.fir@89358.4]
  wire  _T_91; // @[MSHR.scala 187:83:chipyard.TestHarness.RocketConfig.fir@89359.4]
  wire  _T_93; // @[MSHR.scala 189:49:chipyard.TestHarness.RocketConfig.fir@89363.4]
  wire  _T_94; // @[MSHR.scala 189:77:chipyard.TestHarness.RocketConfig.fir@89364.4]
  wire  _T_95; // @[MSHR.scala 189:105:chipyard.TestHarness.RocketConfig.fir@89365.4]
  wire  _T_96; // @[MSHR.scala 190:49:chipyard.TestHarness.RocketConfig.fir@89366.4]
  wire  _T_97; // @[MSHR.scala 190:77:chipyard.TestHarness.RocketConfig.fir@89367.4]
  wire  _GEN_7; // @[MSHR.scala 196:35:chipyard.TestHarness.RocketConfig.fir@89372.6]
  wire  _T_99; // @[MSHR.scala 198:21:chipyard.TestHarness.RocketConfig.fir@89376.6]
  wire  _GEN_8; // @[MSHR.scala 198:35:chipyard.TestHarness.RocketConfig.fir@89377.6]
  wire  _GEN_9; // @[MSHR.scala 199:35:chipyard.TestHarness.RocketConfig.fir@89380.6]
  wire  _GEN_11; // @[MSHR.scala 201:35:chipyard.TestHarness.RocketConfig.fir@89386.6]
  wire  _T_100; // @[MSHR.scala 202:23:chipyard.TestHarness.RocketConfig.fir@89389.6]
  wire  _GEN_12; // @[MSHR.scala 202:35:chipyard.TestHarness.RocketConfig.fir@89390.6]
  wire  _GEN_13; // @[MSHR.scala 203:35:chipyard.TestHarness.RocketConfig.fir@89393.6]
  wire  _GEN_14; // @[MSHR.scala 205:20:chipyard.TestHarness.RocketConfig.fir@89396.6]
  wire  _GEN_15; // @[MSHR.scala 205:20:chipyard.TestHarness.RocketConfig.fir@89396.6]
  wire  _GEN_16; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  wire  _GEN_17; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  wire  _GEN_18; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  wire  _GEN_19; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  wire  _GEN_20; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  wire  _GEN_22; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  wire  _GEN_23; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  wire  _GEN_24; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  wire  _GEN_25; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  wire  _GEN_26; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  wire  req_clientBit; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@89404.4]
  wire  _T_102; // @[Parameters.scala 265:5:chipyard.TestHarness.RocketConfig.fir@89406.4]
  wire  _T_103; // @[Parameters.scala 266:13:chipyard.TestHarness.RocketConfig.fir@89407.4]
  wire  _T_104; // @[Parameters.scala 266:42:chipyard.TestHarness.RocketConfig.fir@89408.4]
  wire  _T_105; // @[Parameters.scala 266:33:chipyard.TestHarness.RocketConfig.fir@89409.4]
  wire  _T_106; // @[Parameters.scala 265:16:chipyard.TestHarness.RocketConfig.fir@89410.4]
  wire  _T_107; // @[Parameters.scala 267:14:chipyard.TestHarness.RocketConfig.fir@89411.4]
  wire  _T_108; // @[Parameters.scala 267:52:chipyard.TestHarness.RocketConfig.fir@89412.4]
  wire  _T_109; // @[Parameters.scala 267:42:chipyard.TestHarness.RocketConfig.fir@89413.4]
  wire  _T_110; // @[Parameters.scala 267:89:chipyard.TestHarness.RocketConfig.fir@89414.4]
  wire  _T_111; // @[Parameters.scala 267:80:chipyard.TestHarness.RocketConfig.fir@89415.4]
  wire  req_needT; // @[Parameters.scala 266:70:chipyard.TestHarness.RocketConfig.fir@89416.4]
  wire  _T_116; // @[MSHR.scala 218:67:chipyard.TestHarness.RocketConfig.fir@89423.4]
  wire  _T_117; // @[MSHR.scala 218:40:chipyard.TestHarness.RocketConfig.fir@89424.4]
  wire  req_promoteT; // @[MSHR.scala 218:34:chipyard.TestHarness.RocketConfig.fir@89425.4]
  wire  _T_120; // @[MSHR.scala 221:48:chipyard.TestHarness.RocketConfig.fir@89429.6]
  wire  _T_121; // @[MSHR.scala 222:55:chipyard.TestHarness.RocketConfig.fir@89431.6]
  wire  _T_123; // @[MSHR.scala 222:64:chipyard.TestHarness.RocketConfig.fir@89433.6]
  wire [1:0] _T_124; // @[MSHR.scala 222:40:chipyard.TestHarness.RocketConfig.fir@89434.6]
  wire  _T_126; // @[Parameters.scala 278:43:chipyard.TestHarness.RocketConfig.fir@89437.6]
  wire  _T_127; // @[Parameters.scala 278:34:chipyard.TestHarness.RocketConfig.fir@89438.6]
  wire  _T_128; // @[Parameters.scala 278:75:chipyard.TestHarness.RocketConfig.fir@89439.6]
  wire  _T_129; // @[Parameters.scala 278:66:chipyard.TestHarness.RocketConfig.fir@89440.6]
  wire  _T_130; // @[MSHR.scala 223:56:chipyard.TestHarness.RocketConfig.fir@89441.6]
  wire  _T_131; // @[MSHR.scala 223:52:chipyard.TestHarness.RocketConfig.fir@89442.6]
  wire  _T_132; // @[MSHR.scala 223:50:chipyard.TestHarness.RocketConfig.fir@89443.6]
  wire  _T_134; // @[MSHR.scala 229:54:chipyard.TestHarness.RocketConfig.fir@89453.10]
  wire  _T_135; // @[MSHR.scala 229:52:chipyard.TestHarness.RocketConfig.fir@89454.10]
  wire  _GEN_27; // @[MSHR.scala 226:21:chipyard.TestHarness.RocketConfig.fir@89450.8]
  wire [1:0] _GEN_28; // @[MSHR.scala 226:21:chipyard.TestHarness.RocketConfig.fir@89450.8]
  wire  _GEN_29; // @[MSHR.scala 226:21:chipyard.TestHarness.RocketConfig.fir@89450.8]
  wire  _T_136; // @[MSHR.scala 233:45:chipyard.TestHarness.RocketConfig.fir@89460.8]
  wire  _T_139; // @[MSHR.scala 233:60:chipyard.TestHarness.RocketConfig.fir@89463.8]
  wire [1:0] _T_140; // @[MSHR.scala 235:40:chipyard.TestHarness.RocketConfig.fir@89465.8]
  wire  _T_141; // @[MSHR.scala 236:41:chipyard.TestHarness.RocketConfig.fir@89466.8]
  wire [1:0] _T_143; // @[MSHR.scala 236:55:chipyard.TestHarness.RocketConfig.fir@89468.8]
  wire  _T_144; // @[MSHR.scala 241:72:chipyard.TestHarness.RocketConfig.fir@89469.8]
  wire [1:0] _T_145; // @[MSHR.scala 241:55:chipyard.TestHarness.RocketConfig.fir@89470.8]
  wire  _T_146; // @[Mux.scala 80:60:chipyard.TestHarness.RocketConfig.fir@89471.8]
  wire  _T_148; // @[Mux.scala 80:60:chipyard.TestHarness.RocketConfig.fir@89473.8]
  wire [1:0] _T_149; // @[Mux.scala 80:57:chipyard.TestHarness.RocketConfig.fir@89474.8]
  wire  _T_150; // @[Mux.scala 80:60:chipyard.TestHarness.RocketConfig.fir@89475.8]
  wire [1:0] _T_151; // @[Mux.scala 80:57:chipyard.TestHarness.RocketConfig.fir@89476.8]
  wire [1:0] _T_152; // @[MSHR.scala 236:40:chipyard.TestHarness.RocketConfig.fir@89477.8]
  wire [1:0] _T_153; // @[MSHR.scala 234:38:chipyard.TestHarness.RocketConfig.fir@89478.8]
  wire  _T_156; // @[MSHR.scala 242:40:chipyard.TestHarness.RocketConfig.fir@89482.8]
  wire  _T_157; // @[MSHR.scala 243:40:chipyard.TestHarness.RocketConfig.fir@89483.8]
  wire  _T_158; // @[MSHR.scala 242:88:chipyard.TestHarness.RocketConfig.fir@89484.8]
  wire  _GEN_30; // @[MSHR.scala 225:57:chipyard.TestHarness.RocketConfig.fir@89449.6]
  wire [1:0] _GEN_31; // @[MSHR.scala 225:57:chipyard.TestHarness.RocketConfig.fir@89449.6]
  wire  _GEN_32; // @[MSHR.scala 225:57:chipyard.TestHarness.RocketConfig.fir@89449.6]
  wire  _GEN_33; // @[MSHR.scala 225:57:chipyard.TestHarness.RocketConfig.fir@89449.6]
  wire [11:0] _GEN_34; // @[MSHR.scala 225:57:chipyard.TestHarness.RocketConfig.fir@89449.6]
  wire  _GEN_35; // @[MSHR.scala 220:54:chipyard.TestHarness.RocketConfig.fir@89427.4]
  wire [1:0] _GEN_36; // @[MSHR.scala 220:54:chipyard.TestHarness.RocketConfig.fir@89427.4]
  wire  _GEN_37; // @[MSHR.scala 220:54:chipyard.TestHarness.RocketConfig.fir@89427.4]
  wire  _GEN_38; // @[MSHR.scala 220:54:chipyard.TestHarness.RocketConfig.fir@89427.4]
  wire [11:0] final_meta_writeback_tag; // @[MSHR.scala 220:54:chipyard.TestHarness.RocketConfig.fir@89427.4]
  wire  _T_161; // @[MSHR.scala 251:27:chipyard.TestHarness.RocketConfig.fir@89493.8]
  wire  _T_163; // @[MSHR.scala 251:14:chipyard.TestHarness.RocketConfig.fir@89495.8]
  wire  _T_164; // @[MSHR.scala 251:14:chipyard.TestHarness.RocketConfig.fir@89496.8]
  wire [1:0] _GEN_42; // @[MSHR.scala 249:21:chipyard.TestHarness.RocketConfig.fir@89490.6]
  wire  final_meta_writeback_hit; // @[MSHR.scala 248:20:chipyard.TestHarness.RocketConfig.fir@89489.4]
  wire  final_meta_writeback_dirty; // @[MSHR.scala 248:20:chipyard.TestHarness.RocketConfig.fir@89489.4]
  wire [1:0] final_meta_writeback_state; // @[MSHR.scala 248:20:chipyard.TestHarness.RocketConfig.fir@89489.4]
  wire  final_meta_writeback_clients; // @[MSHR.scala 248:20:chipyard.TestHarness.RocketConfig.fir@89489.4]
  wire  _T_167; // @[MSHR.scala 273:47:chipyard.TestHarness.RocketConfig.fir@89521.4]
  wire  _T_168; // @[MSHR.scala 273:64:chipyard.TestHarness.RocketConfig.fir@89522.4]
  wire  honour_BtoT; // @[MSHR.scala 273:30:chipyard.TestHarness.RocketConfig.fir@89523.4]
  wire  _T_169; // @[MSHR.scala 276:38:chipyard.TestHarness.RocketConfig.fir@89524.4]
  wire  _T_173; // @[Parameters.scala 275:87:chipyard.TestHarness.RocketConfig.fir@89528.4]
  wire  _T_174; // @[Parameters.scala 275:77:chipyard.TestHarness.RocketConfig.fir@89529.4]
  wire  _T_175; // @[MSHR.scala 276:57:chipyard.TestHarness.RocketConfig.fir@89530.4]
  wire  excluded_client; // @[MSHR.scala 276:28:chipyard.TestHarness.RocketConfig.fir@89531.4]
  wire [1:0] _T_176; // @[MSHR.scala 279:56:chipyard.TestHarness.RocketConfig.fir@89534.4]
  wire [1:0] _T_177; // @[MSHR.scala 279:41:chipyard.TestHarness.RocketConfig.fir@89535.4]
  wire  _T_178; // @[MSHR.scala 280:51:chipyard.TestHarness.RocketConfig.fir@89537.4]
  wire  _T_179; // @[MSHR.scala 281:55:chipyard.TestHarness.RocketConfig.fir@89538.4]
  wire  _T_181; // @[MSHR.scala 281:71:chipyard.TestHarness.RocketConfig.fir@89540.4]
  wire  _T_182; // @[MSHR.scala 281:38:chipyard.TestHarness.RocketConfig.fir@89541.4]
  wire [1:0] _T_185; // @[MSHR.scala 283:97:chipyard.TestHarness.RocketConfig.fir@89546.4]
  wire [2:0] _T_186; // @[MSHR.scala 283:61:chipyard.TestHarness.RocketConfig.fir@89547.4]
  wire  _T_190; // @[MSHR.scala 286:53:chipyard.TestHarness.RocketConfig.fir@89554.4]
  wire  _T_191; // @[MSHR.scala 286:51:chipyard.TestHarness.RocketConfig.fir@89555.4]
  wire  _T_195; // @[MSHR.scala 295:42:chipyard.TestHarness.RocketConfig.fir@89568.4]
  wire [1:0] _T_197; // @[MSHR.scala 297:53:chipyard.TestHarness.RocketConfig.fir@89571.4]
  wire [1:0] _T_198; // @[MSHR.scala 298:53:chipyard.TestHarness.RocketConfig.fir@89572.4]
  wire  _T_199; // @[Mux.scala 80:60:chipyard.TestHarness.RocketConfig.fir@89573.4]
  wire [2:0] _T_200; // @[Mux.scala 80:57:chipyard.TestHarness.RocketConfig.fir@89574.4]
  wire  _T_201; // @[Mux.scala 80:60:chipyard.TestHarness.RocketConfig.fir@89575.4]
  wire [2:0] _T_202; // @[Mux.scala 80:57:chipyard.TestHarness.RocketConfig.fir@89576.4]
  wire  _T_203; // @[Mux.scala 80:60:chipyard.TestHarness.RocketConfig.fir@89577.4]
  wire [2:0] _T_204; // @[Mux.scala 80:57:chipyard.TestHarness.RocketConfig.fir@89578.4]
  wire  _T_212; // @[MSHR.scala 315:32:chipyard.TestHarness.RocketConfig.fir@89600.6]
  wire [1:0] _T_214; // @[MSHR.scala 316:32:chipyard.TestHarness.RocketConfig.fir@89606.8]
  wire [2:0] _T_216; // @[MSHR.scala 317:39:chipyard.TestHarness.RocketConfig.fir@89612.10]
  wire [2:0] _T_217; // @[MSHR.scala 317:76:chipyard.TestHarness.RocketConfig.fir@89613.10]
  wire [2:0] _T_218; // @[MSHR.scala 317:32:chipyard.TestHarness.RocketConfig.fir@89614.10]
  wire [3:0] _GEN_49; // @[Conditional.scala 39:67:chipyard.TestHarness.RocketConfig.fir@89611.8]
  wire [3:0] _GEN_50; // @[Conditional.scala 39:67:chipyard.TestHarness.RocketConfig.fir@89605.6]
  wire [3:0] _GEN_51; // @[Conditional.scala 40:58:chipyard.TestHarness.RocketConfig.fir@89599.4]
  wire  _T_220; // @[MSHR.scala 320:11:chipyard.TestHarness.RocketConfig.fir@89622.4]
  wire [3:0] evict; // @[MSHR.scala 320:17:chipyard.TestHarness.RocketConfig.fir@89623.4]
  wire [3:0] before_; // @[MSHR.scala 320:17:chipyard.TestHarness.RocketConfig.fir@89654.4]
  wire  _T_232; // @[MSHR.scala 312:27:chipyard.TestHarness.RocketConfig.fir@89659.4]
  wire  _T_233; // @[Conditional.scala 37:30:chipyard.TestHarness.RocketConfig.fir@89660.4]
  wire  _T_234; // @[MSHR.scala 315:32:chipyard.TestHarness.RocketConfig.fir@89662.6]
  wire  _T_235; // @[Conditional.scala 37:30:chipyard.TestHarness.RocketConfig.fir@89666.6]
  wire [1:0] _T_236; // @[MSHR.scala 316:32:chipyard.TestHarness.RocketConfig.fir@89668.8]
  wire  _T_237; // @[Conditional.scala 37:30:chipyard.TestHarness.RocketConfig.fir@89672.8]
  wire [2:0] _T_238; // @[MSHR.scala 317:39:chipyard.TestHarness.RocketConfig.fir@89674.10]
  wire [2:0] _T_239; // @[MSHR.scala 317:76:chipyard.TestHarness.RocketConfig.fir@89675.10]
  wire [2:0] _T_240; // @[MSHR.scala 317:32:chipyard.TestHarness.RocketConfig.fir@89676.10]
  wire [3:0] _GEN_59; // @[Conditional.scala 39:67:chipyard.TestHarness.RocketConfig.fir@89673.8]
  wire [3:0] _GEN_60; // @[Conditional.scala 39:67:chipyard.TestHarness.RocketConfig.fir@89667.6]
  wire [3:0] after; // @[Conditional.scala 40:58:chipyard.TestHarness.RocketConfig.fir@89661.4]
  wire  _T_245; // @[MSHR.scala 360:42:chipyard.TestHarness.RocketConfig.fir@89690.4]
  wire  _T_246; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89692.6]
  wire  _T_247; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89693.6]
  wire  _T_249; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89695.6]
  wire  _T_250; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89696.6]
  wire  _T_251; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89701.6]
  wire  _T_252; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89702.6]
  wire  _T_254; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89704.6]
  wire  _T_255; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89705.6]
  wire  _T_256; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89710.6]
  wire  _T_257; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89711.6]
  wire  _T_259; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89713.6]
  wire  _T_260; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89714.6]
  wire  _T_261; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89719.6]
  wire  _T_262; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89720.6]
  wire  _T_264; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89722.6]
  wire  _T_265; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89723.6]
  wire  _T_267; // @[MSHR.scala 363:13:chipyard.TestHarness.RocketConfig.fir@89729.6]
  wire  _T_269; // @[MSHR.scala 364:13:chipyard.TestHarness.RocketConfig.fir@89731.6]
  wire  _T_271; // @[MSHR.scala 365:13:chipyard.TestHarness.RocketConfig.fir@89733.6]
  wire  _T_273; // @[MSHR.scala 366:13:chipyard.TestHarness.RocketConfig.fir@89735.6]
  wire  _T_275; // @[MSHR.scala 367:13:chipyard.TestHarness.RocketConfig.fir@89737.6]
  wire  _T_277; // @[MSHR.scala 368:13:chipyard.TestHarness.RocketConfig.fir@89739.6]
  wire  _T_280; // @[MSHR.scala 371:35:chipyard.TestHarness.RocketConfig.fir@89743.4]
  wire  _T_281; // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89745.6]
  wire  _T_282; // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89746.6]
  wire  _T_283; // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89747.6]
  wire  _T_284; // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89748.6]
  wire  _T_286; // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89750.6]
  wire  _T_287; // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89751.6]
  wire  _T_289; // @[MSHR.scala 373:15:chipyard.TestHarness.RocketConfig.fir@89757.6]
  wire  _T_290; // @[MSHR.scala 373:15:chipyard.TestHarness.RocketConfig.fir@89758.6]
  wire  _T_291; // @[MSHR.scala 373:15:chipyard.TestHarness.RocketConfig.fir@89759.6]
  wire  _T_293; // @[MSHR.scala 373:15:chipyard.TestHarness.RocketConfig.fir@89761.6]
  wire  _T_294; // @[MSHR.scala 373:15:chipyard.TestHarness.RocketConfig.fir@89762.6]
  wire  _T_296; // @[MSHR.scala 374:15:chipyard.TestHarness.RocketConfig.fir@89768.6]
  wire  _T_299; // @[MSHR.scala 375:15:chipyard.TestHarness.RocketConfig.fir@89771.6]
  wire  _T_300; // @[MSHR.scala 375:15:chipyard.TestHarness.RocketConfig.fir@89772.6]
  wire  _T_301; // @[MSHR.scala 375:15:chipyard.TestHarness.RocketConfig.fir@89773.6]
  wire  _T_303; // @[MSHR.scala 375:15:chipyard.TestHarness.RocketConfig.fir@89775.6]
  wire  _T_304; // @[MSHR.scala 375:15:chipyard.TestHarness.RocketConfig.fir@89776.6]
  wire  _T_306; // @[MSHR.scala 376:15:chipyard.TestHarness.RocketConfig.fir@89782.6]
  wire  _T_307; // @[MSHR.scala 376:15:chipyard.TestHarness.RocketConfig.fir@89783.6]
  wire  _T_308; // @[MSHR.scala 376:15:chipyard.TestHarness.RocketConfig.fir@89784.6]
  wire  _T_310; // @[MSHR.scala 376:15:chipyard.TestHarness.RocketConfig.fir@89786.6]
  wire  _T_311; // @[MSHR.scala 376:15:chipyard.TestHarness.RocketConfig.fir@89787.6]
  wire  _T_313; // @[MSHR.scala 377:15:chipyard.TestHarness.RocketConfig.fir@89793.6]
  wire  _T_316; // @[MSHR.scala 378:15:chipyard.TestHarness.RocketConfig.fir@89796.6]
  wire  _T_319; // @[MSHR.scala 379:15:chipyard.TestHarness.RocketConfig.fir@89799.6]
  wire  _T_320; // @[MSHR.scala 379:15:chipyard.TestHarness.RocketConfig.fir@89800.6]
  wire  _T_321; // @[MSHR.scala 379:15:chipyard.TestHarness.RocketConfig.fir@89801.6]
  wire  _T_323; // @[MSHR.scala 379:15:chipyard.TestHarness.RocketConfig.fir@89803.6]
  wire  _T_324; // @[MSHR.scala 379:15:chipyard.TestHarness.RocketConfig.fir@89804.6]
  wire  _T_326; // @[MSHR.scala 381:15:chipyard.TestHarness.RocketConfig.fir@89810.6]
  wire  _T_327; // @[MSHR.scala 381:15:chipyard.TestHarness.RocketConfig.fir@89811.6]
  wire  _T_328; // @[MSHR.scala 381:15:chipyard.TestHarness.RocketConfig.fir@89812.6]
  wire  _T_330; // @[MSHR.scala 381:15:chipyard.TestHarness.RocketConfig.fir@89814.6]
  wire  _T_331; // @[MSHR.scala 381:15:chipyard.TestHarness.RocketConfig.fir@89815.6]
  wire  _T_334; // @[MSHR.scala 382:15:chipyard.TestHarness.RocketConfig.fir@89822.6]
  wire  _T_335; // @[MSHR.scala 382:15:chipyard.TestHarness.RocketConfig.fir@89823.6]
  wire  _T_337; // @[MSHR.scala 382:15:chipyard.TestHarness.RocketConfig.fir@89825.6]
  wire  _T_338; // @[MSHR.scala 382:15:chipyard.TestHarness.RocketConfig.fir@89826.6]
  wire  _T_341; // @[MSHR.scala 383:15:chipyard.TestHarness.RocketConfig.fir@89833.6]
  wire  _T_342; // @[MSHR.scala 383:15:chipyard.TestHarness.RocketConfig.fir@89834.6]
  wire  _T_344; // @[MSHR.scala 383:15:chipyard.TestHarness.RocketConfig.fir@89836.6]
  wire  _T_345; // @[MSHR.scala 383:15:chipyard.TestHarness.RocketConfig.fir@89837.6]
  wire  _T_348; // @[MSHR.scala 384:15:chipyard.TestHarness.RocketConfig.fir@89844.6]
  wire  _T_349; // @[MSHR.scala 384:15:chipyard.TestHarness.RocketConfig.fir@89845.6]
  wire  _T_351; // @[MSHR.scala 384:15:chipyard.TestHarness.RocketConfig.fir@89847.6]
  wire  _T_352; // @[MSHR.scala 384:15:chipyard.TestHarness.RocketConfig.fir@89848.6]
  wire  _T_355; // @[MSHR.scala 385:15:chipyard.TestHarness.RocketConfig.fir@89855.6]
  wire  _T_356; // @[MSHR.scala 385:15:chipyard.TestHarness.RocketConfig.fir@89856.6]
  wire  _T_358; // @[MSHR.scala 385:15:chipyard.TestHarness.RocketConfig.fir@89858.6]
  wire  _T_359; // @[MSHR.scala 385:15:chipyard.TestHarness.RocketConfig.fir@89859.6]
  wire  _T_362; // @[MSHR.scala 386:15:chipyard.TestHarness.RocketConfig.fir@89866.6]
  wire  _T_363; // @[MSHR.scala 386:15:chipyard.TestHarness.RocketConfig.fir@89867.6]
  wire  _T_365; // @[MSHR.scala 386:15:chipyard.TestHarness.RocketConfig.fir@89869.6]
  wire  _T_366; // @[MSHR.scala 386:15:chipyard.TestHarness.RocketConfig.fir@89870.6]
  wire  _T_369; // @[MSHR.scala 387:15:chipyard.TestHarness.RocketConfig.fir@89877.6]
  wire  _T_370; // @[MSHR.scala 387:15:chipyard.TestHarness.RocketConfig.fir@89878.6]
  wire  _T_372; // @[MSHR.scala 387:15:chipyard.TestHarness.RocketConfig.fir@89880.6]
  wire  _T_373; // @[MSHR.scala 387:15:chipyard.TestHarness.RocketConfig.fir@89881.6]
  wire  _T_376; // @[MSHR.scala 388:15:chipyard.TestHarness.RocketConfig.fir@89888.6]
  wire  _T_377; // @[MSHR.scala 388:15:chipyard.TestHarness.RocketConfig.fir@89889.6]
  wire  _T_379; // @[MSHR.scala 388:15:chipyard.TestHarness.RocketConfig.fir@89891.6]
  wire  _T_380; // @[MSHR.scala 388:15:chipyard.TestHarness.RocketConfig.fir@89892.6]
  wire  _T_383; // @[MSHR.scala 390:15:chipyard.TestHarness.RocketConfig.fir@89899.6]
  wire  _T_384; // @[MSHR.scala 390:15:chipyard.TestHarness.RocketConfig.fir@89900.6]
  wire  _T_386; // @[MSHR.scala 390:15:chipyard.TestHarness.RocketConfig.fir@89902.6]
  wire  _T_387; // @[MSHR.scala 390:15:chipyard.TestHarness.RocketConfig.fir@89903.6]
  wire  _T_390; // @[MSHR.scala 391:15:chipyard.TestHarness.RocketConfig.fir@89910.6]
  wire  _T_391; // @[MSHR.scala 391:15:chipyard.TestHarness.RocketConfig.fir@89911.6]
  wire  _T_393; // @[MSHR.scala 391:15:chipyard.TestHarness.RocketConfig.fir@89913.6]
  wire  _T_394; // @[MSHR.scala 391:15:chipyard.TestHarness.RocketConfig.fir@89914.6]
  wire  _T_397; // @[MSHR.scala 392:15:chipyard.TestHarness.RocketConfig.fir@89921.6]
  wire  _T_398; // @[MSHR.scala 392:15:chipyard.TestHarness.RocketConfig.fir@89922.6]
  wire  _T_400; // @[MSHR.scala 392:15:chipyard.TestHarness.RocketConfig.fir@89924.6]
  wire  _T_401; // @[MSHR.scala 392:15:chipyard.TestHarness.RocketConfig.fir@89925.6]
  wire  _T_404; // @[MSHR.scala 393:15:chipyard.TestHarness.RocketConfig.fir@89932.6]
  wire  _T_405; // @[MSHR.scala 393:15:chipyard.TestHarness.RocketConfig.fir@89933.6]
  wire  _T_407; // @[MSHR.scala 393:15:chipyard.TestHarness.RocketConfig.fir@89935.6]
  wire  _T_408; // @[MSHR.scala 393:15:chipyard.TestHarness.RocketConfig.fir@89936.6]
  wire  _T_411; // @[MSHR.scala 394:15:chipyard.TestHarness.RocketConfig.fir@89943.6]
  wire  _T_412; // @[MSHR.scala 394:15:chipyard.TestHarness.RocketConfig.fir@89944.6]
  wire  _T_414; // @[MSHR.scala 394:15:chipyard.TestHarness.RocketConfig.fir@89946.6]
  wire  _T_415; // @[MSHR.scala 394:15:chipyard.TestHarness.RocketConfig.fir@89947.6]
  wire  _T_418; // @[MSHR.scala 395:15:chipyard.TestHarness.RocketConfig.fir@89954.6]
  wire  _T_419; // @[MSHR.scala 395:15:chipyard.TestHarness.RocketConfig.fir@89955.6]
  wire  _T_421; // @[MSHR.scala 395:15:chipyard.TestHarness.RocketConfig.fir@89957.6]
  wire  _T_422; // @[MSHR.scala 395:15:chipyard.TestHarness.RocketConfig.fir@89958.6]
  wire  _T_425; // @[MSHR.scala 396:15:chipyard.TestHarness.RocketConfig.fir@89965.6]
  wire  _T_426; // @[MSHR.scala 396:15:chipyard.TestHarness.RocketConfig.fir@89966.6]
  wire  _T_428; // @[MSHR.scala 396:15:chipyard.TestHarness.RocketConfig.fir@89968.6]
  wire  _T_429; // @[MSHR.scala 396:15:chipyard.TestHarness.RocketConfig.fir@89969.6]
  wire  _T_432; // @[MSHR.scala 397:15:chipyard.TestHarness.RocketConfig.fir@89976.6]
  wire  _T_433; // @[MSHR.scala 397:15:chipyard.TestHarness.RocketConfig.fir@89977.6]
  wire  _T_435; // @[MSHR.scala 397:15:chipyard.TestHarness.RocketConfig.fir@89979.6]
  wire  _T_436; // @[MSHR.scala 397:15:chipyard.TestHarness.RocketConfig.fir@89980.6]
  wire  _T_439; // @[MSHR.scala 399:15:chipyard.TestHarness.RocketConfig.fir@89987.6]
  wire  _T_440; // @[MSHR.scala 399:15:chipyard.TestHarness.RocketConfig.fir@89988.6]
  wire  _T_442; // @[MSHR.scala 399:15:chipyard.TestHarness.RocketConfig.fir@89990.6]
  wire  _T_443; // @[MSHR.scala 399:15:chipyard.TestHarness.RocketConfig.fir@89991.6]
  wire  _T_446; // @[MSHR.scala 400:15:chipyard.TestHarness.RocketConfig.fir@89998.6]
  wire  _T_447; // @[MSHR.scala 400:15:chipyard.TestHarness.RocketConfig.fir@89999.6]
  wire  _T_449; // @[MSHR.scala 400:15:chipyard.TestHarness.RocketConfig.fir@90001.6]
  wire  _T_450; // @[MSHR.scala 400:15:chipyard.TestHarness.RocketConfig.fir@90002.6]
  wire  _T_453; // @[MSHR.scala 401:15:chipyard.TestHarness.RocketConfig.fir@90009.6]
  wire  _T_454; // @[MSHR.scala 401:15:chipyard.TestHarness.RocketConfig.fir@90010.6]
  wire  _T_456; // @[MSHR.scala 401:15:chipyard.TestHarness.RocketConfig.fir@90012.6]
  wire  _T_457; // @[MSHR.scala 401:15:chipyard.TestHarness.RocketConfig.fir@90013.6]
  wire  _T_460; // @[MSHR.scala 402:15:chipyard.TestHarness.RocketConfig.fir@90020.6]
  wire  _T_461; // @[MSHR.scala 402:15:chipyard.TestHarness.RocketConfig.fir@90021.6]
  wire  _T_463; // @[MSHR.scala 402:15:chipyard.TestHarness.RocketConfig.fir@90023.6]
  wire  _T_464; // @[MSHR.scala 402:15:chipyard.TestHarness.RocketConfig.fir@90024.6]
  wire  _T_470; // @[MSHR.scala 404:15:chipyard.TestHarness.RocketConfig.fir@90034.6]
  wire  _T_471; // @[MSHR.scala 404:15:chipyard.TestHarness.RocketConfig.fir@90035.6]
  wire  _T_473; // @[MSHR.scala 404:15:chipyard.TestHarness.RocketConfig.fir@90037.6]
  wire  _T_474; // @[MSHR.scala 404:15:chipyard.TestHarness.RocketConfig.fir@90038.6]
  wire  _T_480; // @[MSHR.scala 406:15:chipyard.TestHarness.RocketConfig.fir@90048.6]
  wire  _T_481; // @[MSHR.scala 406:15:chipyard.TestHarness.RocketConfig.fir@90049.6]
  wire  _T_483; // @[MSHR.scala 406:15:chipyard.TestHarness.RocketConfig.fir@90051.6]
  wire  _T_484; // @[MSHR.scala 406:15:chipyard.TestHarness.RocketConfig.fir@90052.6]
  wire  _T_487; // @[MSHR.scala 408:15:chipyard.TestHarness.RocketConfig.fir@90059.6]
  wire  _T_488; // @[MSHR.scala 408:15:chipyard.TestHarness.RocketConfig.fir@90060.6]
  wire  _T_490; // @[MSHR.scala 408:15:chipyard.TestHarness.RocketConfig.fir@90062.6]
  wire  _T_491; // @[MSHR.scala 408:15:chipyard.TestHarness.RocketConfig.fir@90063.6]
  wire  _T_494; // @[MSHR.scala 409:15:chipyard.TestHarness.RocketConfig.fir@90070.6]
  wire  _T_495; // @[MSHR.scala 409:15:chipyard.TestHarness.RocketConfig.fir@90071.6]
  wire  _T_497; // @[MSHR.scala 409:15:chipyard.TestHarness.RocketConfig.fir@90073.6]
  wire  _T_498; // @[MSHR.scala 409:15:chipyard.TestHarness.RocketConfig.fir@90074.6]
  wire  _T_501; // @[MSHR.scala 410:15:chipyard.TestHarness.RocketConfig.fir@90081.6]
  wire  _T_502; // @[MSHR.scala 410:15:chipyard.TestHarness.RocketConfig.fir@90082.6]
  wire  _T_504; // @[MSHR.scala 410:15:chipyard.TestHarness.RocketConfig.fir@90084.6]
  wire  _T_505; // @[MSHR.scala 410:15:chipyard.TestHarness.RocketConfig.fir@90085.6]
  wire  _T_514; // @[MSHR.scala 413:15:chipyard.TestHarness.RocketConfig.fir@90098.6]
  wire  _T_515; // @[MSHR.scala 413:15:chipyard.TestHarness.RocketConfig.fir@90099.6]
  wire  _T_517; // @[MSHR.scala 413:15:chipyard.TestHarness.RocketConfig.fir@90101.6]
  wire  _T_518; // @[MSHR.scala 413:15:chipyard.TestHarness.RocketConfig.fir@90102.6]
  wire  _T_524; // @[MSHR.scala 415:15:chipyard.TestHarness.RocketConfig.fir@90112.6]
  wire  _T_525; // @[MSHR.scala 415:15:chipyard.TestHarness.RocketConfig.fir@90113.6]
  wire  _T_527; // @[MSHR.scala 415:15:chipyard.TestHarness.RocketConfig.fir@90115.6]
  wire  _T_528; // @[MSHR.scala 415:15:chipyard.TestHarness.RocketConfig.fir@90116.6]
  wire  _T_531; // @[MSHR.scala 417:15:chipyard.TestHarness.RocketConfig.fir@90123.6]
  wire  _T_532; // @[MSHR.scala 417:15:chipyard.TestHarness.RocketConfig.fir@90124.6]
  wire  _T_534; // @[MSHR.scala 417:15:chipyard.TestHarness.RocketConfig.fir@90126.6]
  wire  _T_535; // @[MSHR.scala 417:15:chipyard.TestHarness.RocketConfig.fir@90127.6]
  wire  _T_538; // @[MSHR.scala 418:15:chipyard.TestHarness.RocketConfig.fir@90134.6]
  wire  _T_539; // @[MSHR.scala 418:15:chipyard.TestHarness.RocketConfig.fir@90135.6]
  wire  _T_541; // @[MSHR.scala 418:15:chipyard.TestHarness.RocketConfig.fir@90137.6]
  wire  _T_542; // @[MSHR.scala 418:15:chipyard.TestHarness.RocketConfig.fir@90138.6]
  wire  _T_545; // @[MSHR.scala 419:15:chipyard.TestHarness.RocketConfig.fir@90145.6]
  wire  _T_546; // @[MSHR.scala 419:15:chipyard.TestHarness.RocketConfig.fir@90146.6]
  wire  _T_548; // @[MSHR.scala 419:15:chipyard.TestHarness.RocketConfig.fir@90148.6]
  wire  _T_549; // @[MSHR.scala 419:15:chipyard.TestHarness.RocketConfig.fir@90149.6]
  wire  _T_552; // @[MSHR.scala 420:15:chipyard.TestHarness.RocketConfig.fir@90156.6]
  wire  _T_553; // @[MSHR.scala 420:15:chipyard.TestHarness.RocketConfig.fir@90157.6]
  wire  _T_555; // @[MSHR.scala 420:15:chipyard.TestHarness.RocketConfig.fir@90159.6]
  wire  _T_556; // @[MSHR.scala 420:15:chipyard.TestHarness.RocketConfig.fir@90160.6]
  wire  _T_559; // @[MSHR.scala 421:15:chipyard.TestHarness.RocketConfig.fir@90167.6]
  wire  _T_560; // @[MSHR.scala 421:15:chipyard.TestHarness.RocketConfig.fir@90168.6]
  wire  _T_562; // @[MSHR.scala 421:15:chipyard.TestHarness.RocketConfig.fir@90170.6]
  wire  _T_563; // @[MSHR.scala 421:15:chipyard.TestHarness.RocketConfig.fir@90171.6]
  wire  _T_566; // @[MSHR.scala 422:15:chipyard.TestHarness.RocketConfig.fir@90178.6]
  wire  _T_567; // @[MSHR.scala 422:15:chipyard.TestHarness.RocketConfig.fir@90179.6]
  wire  _T_569; // @[MSHR.scala 422:15:chipyard.TestHarness.RocketConfig.fir@90181.6]
  wire  _T_570; // @[MSHR.scala 422:15:chipyard.TestHarness.RocketConfig.fir@90182.6]
  wire  _T_573; // @[MSHR.scala 423:15:chipyard.TestHarness.RocketConfig.fir@90189.6]
  wire  _T_574; // @[MSHR.scala 423:15:chipyard.TestHarness.RocketConfig.fir@90190.6]
  wire  _T_576; // @[MSHR.scala 423:15:chipyard.TestHarness.RocketConfig.fir@90192.6]
  wire  _T_577; // @[MSHR.scala 423:15:chipyard.TestHarness.RocketConfig.fir@90193.6]
  wire  _T_583; // @[MSHR.scala 426:15:chipyard.TestHarness.RocketConfig.fir@90203.6]
  wire  _T_584; // @[MSHR.scala 426:15:chipyard.TestHarness.RocketConfig.fir@90204.6]
  wire  _T_586; // @[MSHR.scala 426:15:chipyard.TestHarness.RocketConfig.fir@90206.6]
  wire  _T_587; // @[MSHR.scala 426:15:chipyard.TestHarness.RocketConfig.fir@90207.6]
  wire  _T_590; // @[MSHR.scala 427:15:chipyard.TestHarness.RocketConfig.fir@90214.6]
  wire  _T_591; // @[MSHR.scala 427:15:chipyard.TestHarness.RocketConfig.fir@90215.6]
  wire  _T_593; // @[MSHR.scala 427:15:chipyard.TestHarness.RocketConfig.fir@90217.6]
  wire  _T_594; // @[MSHR.scala 427:15:chipyard.TestHarness.RocketConfig.fir@90218.6]
  wire  _T_597; // @[MSHR.scala 428:15:chipyard.TestHarness.RocketConfig.fir@90225.6]
  wire  _T_598; // @[MSHR.scala 428:15:chipyard.TestHarness.RocketConfig.fir@90226.6]
  wire  _T_600; // @[MSHR.scala 428:15:chipyard.TestHarness.RocketConfig.fir@90228.6]
  wire  _T_601; // @[MSHR.scala 428:15:chipyard.TestHarness.RocketConfig.fir@90229.6]
  wire  _T_604; // @[MSHR.scala 429:15:chipyard.TestHarness.RocketConfig.fir@90236.6]
  wire  _T_605; // @[MSHR.scala 429:15:chipyard.TestHarness.RocketConfig.fir@90237.6]
  wire  _T_607; // @[MSHR.scala 429:15:chipyard.TestHarness.RocketConfig.fir@90239.6]
  wire  _T_608; // @[MSHR.scala 429:15:chipyard.TestHarness.RocketConfig.fir@90240.6]
  wire  _T_611; // @[MSHR.scala 430:15:chipyard.TestHarness.RocketConfig.fir@90247.6]
  wire  _T_612; // @[MSHR.scala 430:15:chipyard.TestHarness.RocketConfig.fir@90248.6]
  wire  _T_614; // @[MSHR.scala 430:15:chipyard.TestHarness.RocketConfig.fir@90250.6]
  wire  _T_615; // @[MSHR.scala 430:15:chipyard.TestHarness.RocketConfig.fir@90251.6]
  wire  _T_621; // @[MSHR.scala 432:15:chipyard.TestHarness.RocketConfig.fir@90261.6]
  wire  _T_622; // @[MSHR.scala 432:15:chipyard.TestHarness.RocketConfig.fir@90262.6]
  wire  _T_624; // @[MSHR.scala 432:15:chipyard.TestHarness.RocketConfig.fir@90264.6]
  wire  _T_625; // @[MSHR.scala 432:15:chipyard.TestHarness.RocketConfig.fir@90265.6]
  wire  _T_631; // @[MSHR.scala 435:15:chipyard.TestHarness.RocketConfig.fir@90275.6]
  wire  _T_632; // @[MSHR.scala 435:15:chipyard.TestHarness.RocketConfig.fir@90276.6]
  wire  _T_634; // @[MSHR.scala 435:15:chipyard.TestHarness.RocketConfig.fir@90278.6]
  wire  _T_635; // @[MSHR.scala 435:15:chipyard.TestHarness.RocketConfig.fir@90279.6]
  wire  _T_638; // @[MSHR.scala 436:15:chipyard.TestHarness.RocketConfig.fir@90286.6]
  wire  _T_639; // @[MSHR.scala 436:15:chipyard.TestHarness.RocketConfig.fir@90287.6]
  wire  _T_641; // @[MSHR.scala 436:15:chipyard.TestHarness.RocketConfig.fir@90289.6]
  wire  _T_642; // @[MSHR.scala 436:15:chipyard.TestHarness.RocketConfig.fir@90290.6]
  wire  _T_645; // @[MSHR.scala 437:15:chipyard.TestHarness.RocketConfig.fir@90297.6]
  wire  _T_646; // @[MSHR.scala 437:15:chipyard.TestHarness.RocketConfig.fir@90298.6]
  wire  _T_648; // @[MSHR.scala 437:15:chipyard.TestHarness.RocketConfig.fir@90300.6]
  wire  _T_649; // @[MSHR.scala 437:15:chipyard.TestHarness.RocketConfig.fir@90301.6]
  wire  _T_667; // @[MSHR.scala 444:15:chipyard.TestHarness.RocketConfig.fir@90323.6]
  wire  _T_668; // @[MSHR.scala 444:15:chipyard.TestHarness.RocketConfig.fir@90324.6]
  wire  _T_670; // @[MSHR.scala 444:15:chipyard.TestHarness.RocketConfig.fir@90326.6]
  wire  _T_671; // @[MSHR.scala 444:15:chipyard.TestHarness.RocketConfig.fir@90327.6]
  wire  _T_674; // @[MSHR.scala 445:15:chipyard.TestHarness.RocketConfig.fir@90334.6]
  wire  _T_675; // @[MSHR.scala 445:15:chipyard.TestHarness.RocketConfig.fir@90335.6]
  wire  _T_677; // @[MSHR.scala 445:15:chipyard.TestHarness.RocketConfig.fir@90337.6]
  wire  _T_678; // @[MSHR.scala 445:15:chipyard.TestHarness.RocketConfig.fir@90338.6]
  wire  _T_681; // @[MSHR.scala 446:15:chipyard.TestHarness.RocketConfig.fir@90345.6]
  wire  _T_682; // @[MSHR.scala 446:15:chipyard.TestHarness.RocketConfig.fir@90346.6]
  wire  _T_684; // @[MSHR.scala 446:15:chipyard.TestHarness.RocketConfig.fir@90348.6]
  wire  _T_685; // @[MSHR.scala 446:15:chipyard.TestHarness.RocketConfig.fir@90349.6]
  wire  _T_688; // @[MSHR.scala 447:15:chipyard.TestHarness.RocketConfig.fir@90356.6]
  wire  _T_689; // @[MSHR.scala 447:15:chipyard.TestHarness.RocketConfig.fir@90357.6]
  wire  _T_691; // @[MSHR.scala 447:15:chipyard.TestHarness.RocketConfig.fir@90359.6]
  wire  _T_692; // @[MSHR.scala 447:15:chipyard.TestHarness.RocketConfig.fir@90360.6]
  wire  _T_695; // @[MSHR.scala 448:15:chipyard.TestHarness.RocketConfig.fir@90367.6]
  wire  _T_696; // @[MSHR.scala 448:15:chipyard.TestHarness.RocketConfig.fir@90368.6]
  wire  _T_698; // @[MSHR.scala 448:15:chipyard.TestHarness.RocketConfig.fir@90370.6]
  wire  _T_699; // @[MSHR.scala 448:15:chipyard.TestHarness.RocketConfig.fir@90371.6]
  wire  _T_708; // @[MSHR.scala 451:15:chipyard.TestHarness.RocketConfig.fir@90384.6]
  wire  _T_709; // @[MSHR.scala 451:15:chipyard.TestHarness.RocketConfig.fir@90385.6]
  wire  _T_711; // @[MSHR.scala 451:15:chipyard.TestHarness.RocketConfig.fir@90387.6]
  wire  _T_712; // @[MSHR.scala 451:15:chipyard.TestHarness.RocketConfig.fir@90388.6]
  wire  probe_bit; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@90394.4]
  wire  _T_713; // @[MSHR.scala 456:33:chipyard.TestHarness.RocketConfig.fir@90395.4]
  wire  last_probe; // @[MSHR.scala 456:46:chipyard.TestHarness.RocketConfig.fir@90398.4]
  wire  _T_716; // @[Parameters.scala 278:11:chipyard.TestHarness.RocketConfig.fir@90399.4]
  wire  _T_717; // @[Parameters.scala 278:43:chipyard.TestHarness.RocketConfig.fir@90400.4]
  wire  _T_718; // @[Parameters.scala 278:34:chipyard.TestHarness.RocketConfig.fir@90401.4]
  wire  _T_719; // @[Parameters.scala 278:75:chipyard.TestHarness.RocketConfig.fir@90402.4]
  wire  probe_toN; // @[Parameters.scala 278:66:chipyard.TestHarness.RocketConfig.fir@90403.4]
  wire  _T_726; // @[MSHR.scala 465:35:chipyard.TestHarness.RocketConfig.fir@90412.6]
  wire  _T_727; // @[MSHR.scala 465:30:chipyard.TestHarness.RocketConfig.fir@90413.6]
  wire  _T_730; // @[MSHR.scala 467:42:chipyard.TestHarness.RocketConfig.fir@90418.6]
  wire  _T_731; // @[MSHR.scala 468:55:chipyard.TestHarness.RocketConfig.fir@90420.6]
  wire  _T_732; // @[MSHR.scala 468:40:chipyard.TestHarness.RocketConfig.fir@90421.6]
  wire  _T_733; // @[MSHR.scala 469:42:chipyard.TestHarness.RocketConfig.fir@90423.6]
  wire  _T_735; // @[MSHR.scala 470:40:chipyard.TestHarness.RocketConfig.fir@90426.6]
  wire  _T_736; // @[MSHR.scala 472:77:chipyard.TestHarness.RocketConfig.fir@90428.6]
  wire  _T_737; // @[MSHR.scala 472:59:chipyard.TestHarness.RocketConfig.fir@90429.6]
  wire  _T_738; // @[MSHR.scala 472:36:chipyard.TestHarness.RocketConfig.fir@90430.6]
  wire  _T_739; // @[MSHR.scala 473:32:chipyard.TestHarness.RocketConfig.fir@90431.6]
  wire  _T_744; // @[MSHR.scala 477:55:chipyard.TestHarness.RocketConfig.fir@90437.6]
  wire  _T_745; // @[MSHR.scala 477:34:chipyard.TestHarness.RocketConfig.fir@90438.6]
  wire  _T_746; // @[MSHR.scala 477:68:chipyard.TestHarness.RocketConfig.fir@90439.6]
  wire  _GEN_63; // @[MSHR.scala 477:91:chipyard.TestHarness.RocketConfig.fir@90440.6]
  wire  _GEN_67; // @[MSHR.scala 458:49:chipyard.TestHarness.RocketConfig.fir@90404.4]
  wire  _GEN_68; // @[MSHR.scala 458:49:chipyard.TestHarness.RocketConfig.fir@90404.4]
  wire  _GEN_69; // @[MSHR.scala 458:49:chipyard.TestHarness.RocketConfig.fir@90404.4]
  wire  _GEN_70; // @[MSHR.scala 458:49:chipyard.TestHarness.RocketConfig.fir@90404.4]
  wire  _GEN_71; // @[MSHR.scala 458:49:chipyard.TestHarness.RocketConfig.fir@90404.4]
  wire  _T_747; // @[MSHR.scala 480:32:chipyard.TestHarness.RocketConfig.fir@90445.6]
  wire  _T_748; // @[MSHR.scala 480:66:chipyard.TestHarness.RocketConfig.fir@90446.6]
  wire  _T_749; // @[MSHR.scala 480:42:chipyard.TestHarness.RocketConfig.fir@90447.6]
  wire  _T_751; // @[MSHR.scala 487:45:chipyard.TestHarness.RocketConfig.fir@90454.8]
  wire  _T_758; // @[MSHR.scala 490:35:chipyard.TestHarness.RocketConfig.fir@90462.8]
  wire  _T_759; // @[MSHR.scala 492:37:chipyard.TestHarness.RocketConfig.fir@90466.8]
  wire  _GEN_73; // @[MSHR.scala 492:53:chipyard.TestHarness.RocketConfig.fir@90467.8]
  wire  _GEN_75; // @[MSHR.scala 480:81:chipyard.TestHarness.RocketConfig.fir@90448.6]
  wire  _GEN_76; // @[MSHR.scala 480:81:chipyard.TestHarness.RocketConfig.fir@90448.6]
  wire  _GEN_78; // @[MSHR.scala 480:81:chipyard.TestHarness.RocketConfig.fir@90448.6]
  wire  _GEN_80; // @[MSHR.scala 480:81:chipyard.TestHarness.RocketConfig.fir@90448.6]
  wire  _GEN_82; // @[MSHR.scala 479:25:chipyard.TestHarness.RocketConfig.fir@90444.4]
  wire  _GEN_83; // @[MSHR.scala 479:25:chipyard.TestHarness.RocketConfig.fir@90444.4]
  wire  _GEN_85; // @[MSHR.scala 479:25:chipyard.TestHarness.RocketConfig.fir@90444.4]
  wire  _GEN_87; // @[MSHR.scala 479:25:chipyard.TestHarness.RocketConfig.fir@90444.4]
  wire  _GEN_88; // @[MSHR.scala 496:25:chipyard.TestHarness.RocketConfig.fir@90471.4]
  wire  _T_760; // @[MSHR.scala 502:40:chipyard.TestHarness.RocketConfig.fir@90477.4]
  wire  new_meta_dirty; // @[MSHR.scala 502:21:chipyard.TestHarness.RocketConfig.fir@90478.4]
  wire [1:0] new_meta_state; // @[MSHR.scala 502:21:chipyard.TestHarness.RocketConfig.fir@90478.4]
  wire  new_meta_clients; // @[MSHR.scala 502:21:chipyard.TestHarness.RocketConfig.fir@90478.4]
  wire  new_meta_hit; // @[MSHR.scala 502:21:chipyard.TestHarness.RocketConfig.fir@90478.4]
  wire  new_request_prio_2; // @[MSHR.scala 503:24:chipyard.TestHarness.RocketConfig.fir@90479.4]
  wire  new_request_control; // @[MSHR.scala 503:24:chipyard.TestHarness.RocketConfig.fir@90479.4]
  wire [2:0] new_request_opcode; // @[MSHR.scala 503:24:chipyard.TestHarness.RocketConfig.fir@90479.4]
  wire [2:0] new_request_param; // @[MSHR.scala 503:24:chipyard.TestHarness.RocketConfig.fir@90479.4]
  wire [2:0] new_request_source; // @[MSHR.scala 503:24:chipyard.TestHarness.RocketConfig.fir@90479.4]
  wire  _T_762; // @[Parameters.scala 265:5:chipyard.TestHarness.RocketConfig.fir@90481.4]
  wire  _T_763; // @[Parameters.scala 266:13:chipyard.TestHarness.RocketConfig.fir@90482.4]
  wire  _T_764; // @[Parameters.scala 266:42:chipyard.TestHarness.RocketConfig.fir@90483.4]
  wire  _T_765; // @[Parameters.scala 266:33:chipyard.TestHarness.RocketConfig.fir@90484.4]
  wire  _T_766; // @[Parameters.scala 265:16:chipyard.TestHarness.RocketConfig.fir@90485.4]
  wire  _T_767; // @[Parameters.scala 267:14:chipyard.TestHarness.RocketConfig.fir@90486.4]
  wire  _T_768; // @[Parameters.scala 267:52:chipyard.TestHarness.RocketConfig.fir@90487.4]
  wire  _T_769; // @[Parameters.scala 267:42:chipyard.TestHarness.RocketConfig.fir@90488.4]
  wire  _T_770; // @[Parameters.scala 267:89:chipyard.TestHarness.RocketConfig.fir@90489.4]
  wire  _T_771; // @[Parameters.scala 267:80:chipyard.TestHarness.RocketConfig.fir@90490.4]
  wire  new_needT; // @[Parameters.scala 266:70:chipyard.TestHarness.RocketConfig.fir@90491.4]
  wire  new_clientBit; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@90492.4]
  wire  _T_775; // @[Parameters.scala 275:87:chipyard.TestHarness.RocketConfig.fir@90496.4]
  wire  _T_776; // @[Parameters.scala 275:77:chipyard.TestHarness.RocketConfig.fir@90497.4]
  wire  new_skipProbe; // @[MSHR.scala 506:26:chipyard.TestHarness.RocketConfig.fir@90498.4]
  wire  _T_791; // @[MSHR.scala 519:11:chipyard.TestHarness.RocketConfig.fir@90534.6]
  wire  _T_793; // @[MSHR.scala 519:11:chipyard.TestHarness.RocketConfig.fir@90536.6]
  wire  _T_794; // @[MSHR.scala 519:11:chipyard.TestHarness.RocketConfig.fir@90537.6]
  wire  _T_796; // @[MSHR.scala 520:11:chipyard.TestHarness.RocketConfig.fir@90543.6]
  wire  _T_798; // @[MSHR.scala 520:11:chipyard.TestHarness.RocketConfig.fir@90545.6]
  wire  _T_799; // @[MSHR.scala 520:11:chipyard.TestHarness.RocketConfig.fir@90546.6]
  wire  _T_806; // @[MSHR.scala 530:13:chipyard.TestHarness.RocketConfig.fir@90559.6]
  wire  _T_807; // @[Decoupled.scala 40:37:chipyard.TestHarness.RocketConfig.fir@90560.6]
  wire  _T_808; // @[MSHR.scala 530:40:chipyard.TestHarness.RocketConfig.fir@90561.6]
  wire  _T_809; // @[MSHR.scala 530:28:chipyard.TestHarness.RocketConfig.fir@90562.6]
  wire  _T_811; // @[MSHR.scala 530:12:chipyard.TestHarness.RocketConfig.fir@90564.6]
  wire  _T_812; // @[MSHR.scala 530:12:chipyard.TestHarness.RocketConfig.fir@90565.6]
  wire  _GEN_94; // @[MSHR.scala 529:28:chipyard.TestHarness.RocketConfig.fir@90558.4]
  wire  _T_814; // @[MSHR.scala 536:28:chipyard.TestHarness.RocketConfig.fir@90574.4]
  wire  _T_817; // @[MSHR.scala 571:38:chipyard.TestHarness.RocketConfig.fir@90606.8]
  wire  _T_818; // @[MSHR.scala 571:35:chipyard.TestHarness.RocketConfig.fir@90607.8]
  wire  _GEN_107; // @[MSHR.scala 571:55:chipyard.TestHarness.RocketConfig.fir@90608.8]
  wire  _T_819; // @[Parameters.scala 281:11:chipyard.TestHarness.RocketConfig.fir@90611.8]
  wire  _T_820; // @[Parameters.scala 281:43:chipyard.TestHarness.RocketConfig.fir@90612.8]
  wire  _T_821; // @[Parameters.scala 281:34:chipyard.TestHarness.RocketConfig.fir@90613.8]
  wire  _T_822; // @[MSHR.scala 575:56:chipyard.TestHarness.RocketConfig.fir@90614.8]
  wire  _T_823; // @[MSHR.scala 575:38:chipyard.TestHarness.RocketConfig.fir@90615.8]
  wire  _GEN_108; // @[MSHR.scala 575:67:chipyard.TestHarness.RocketConfig.fir@90616.8]
  wire  _T_825; // @[Parameters.scala 278:43:chipyard.TestHarness.RocketConfig.fir@90620.8]
  wire  _T_826; // @[Parameters.scala 278:34:chipyard.TestHarness.RocketConfig.fir@90621.8]
  wire  _T_827; // @[Parameters.scala 278:75:chipyard.TestHarness.RocketConfig.fir@90622.8]
  wire  _T_828; // @[Parameters.scala 278:66:chipyard.TestHarness.RocketConfig.fir@90623.8]
  wire  _T_829; // @[MSHR.scala 579:59:chipyard.TestHarness.RocketConfig.fir@90624.8]
  wire  _T_831; // @[MSHR.scala 579:38:chipyard.TestHarness.RocketConfig.fir@90626.8]
  wire  _GEN_109; // @[MSHR.scala 579:89:chipyard.TestHarness.RocketConfig.fir@90627.8]
  wire  _T_833; // @[MSHR.scala 582:14:chipyard.TestHarness.RocketConfig.fir@90631.8]
  wire  _T_834; // @[MSHR.scala 582:14:chipyard.TestHarness.RocketConfig.fir@90632.8]
  wire  _GEN_110; // @[MSHR.scala 592:75:chipyard.TestHarness.RocketConfig.fir@90647.12]
  wire  _GEN_111; // @[MSHR.scala 588:27:chipyard.TestHarness.RocketConfig.fir@90642.10]
  wire  _GEN_112; // @[MSHR.scala 588:27:chipyard.TestHarness.RocketConfig.fir@90642.10]
  wire  _T_838; // @[MSHR.scala 603:13:chipyard.TestHarness.RocketConfig.fir@90656.10]
  wire  _T_839; // @[MSHR.scala 603:45:chipyard.TestHarness.RocketConfig.fir@90657.10]
  wire  _T_840; // @[MSHR.scala 603:27:chipyard.TestHarness.RocketConfig.fir@90658.10]
  wire  _GEN_114; // @[MSHR.scala 603:58:chipyard.TestHarness.RocketConfig.fir@90659.10]
  wire  _GEN_115; // @[MSHR.scala 603:58:chipyard.TestHarness.RocketConfig.fir@90659.10]
  wire  _T_844; // @[MSHR.scala 614:46:chipyard.TestHarness.RocketConfig.fir@90671.10]
  wire  _T_845; // @[MSHR.scala 614:57:chipyard.TestHarness.RocketConfig.fir@90672.10]
  wire  _T_846; // @[MSHR.scala 614:27:chipyard.TestHarness.RocketConfig.fir@90673.10]
  wire  _GEN_116; // @[MSHR.scala 614:72:chipyard.TestHarness.RocketConfig.fir@90674.10]
  wire  _T_848; // @[MSHR.scala 624:24:chipyard.TestHarness.RocketConfig.fir@90683.10]
  wire  _T_849; // @[MSHR.scala 623:55:chipyard.TestHarness.RocketConfig.fir@90684.10]
  wire  _T_850; // @[MSHR.scala 625:33:chipyard.TestHarness.RocketConfig.fir@90685.10]
  wire  _T_851; // @[MSHR.scala 625:31:chipyard.TestHarness.RocketConfig.fir@90686.10]
  wire  _T_853; // @[MSHR.scala 624:53:chipyard.TestHarness.RocketConfig.fir@90688.10]
  wire  _GEN_117; // @[MSHR.scala 625:63:chipyard.TestHarness.RocketConfig.fir@90690.10]
  wire  _GEN_118; // @[MSHR.scala 625:63:chipyard.TestHarness.RocketConfig.fir@90690.10]
  wire  _GEN_119; // @[MSHR.scala 633:88:chipyard.TestHarness.RocketConfig.fir@90700.10]
  wire  _GEN_120; // @[MSHR.scala 633:88:chipyard.TestHarness.RocketConfig.fir@90700.10]
  wire  _T_860; // @[MSHR.scala 638:36:chipyard.TestHarness.RocketConfig.fir@90706.10]
  wire  _T_862; // @[MSHR.scala 638:52:chipyard.TestHarness.RocketConfig.fir@90708.10]
  wire  _GEN_121; // @[MSHR.scala 638:72:chipyard.TestHarness.RocketConfig.fir@90709.10]
  wire  _GEN_122; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  wire  _GEN_123; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  wire  _GEN_124; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  wire  _GEN_126; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  wire  _GEN_127; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  wire  _GEN_128; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  wire  _GEN_129; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  wire  _GEN_130; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  wire  _GEN_131; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  wire  _GEN_132; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  wire  _GEN_133; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  wire  _GEN_134; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  wire  _GEN_135; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  wire  _GEN_136; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  wire  _GEN_137; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  wire  _GEN_138; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_150; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_151; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_152; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_153; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_154; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_155; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_156; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_157; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_158; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_159; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_160; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_161; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_162; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_163; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_165; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_166; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_167; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_168; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  wire  _GEN_170; // @[MSHR.scala 102:14:chipyard.TestHarness.RocketConfig.fir@89185.10]
  wire  _GEN_174; // @[MSHR.scala 106:14:chipyard.TestHarness.RocketConfig.fir@89204.10]
  wire  _GEN_176; // @[MSHR.scala 109:14:chipyard.TestHarness.RocketConfig.fir@89215.10]
  wire  _GEN_180; // @[MSHR.scala 251:14:chipyard.TestHarness.RocketConfig.fir@89498.10]
  wire  _GEN_182; // @[MSHR.scala 582:14:chipyard.TestHarness.RocketConfig.fir@90634.10]
  assign _T = meta_state == 2'h0; // @[MSHR.scala 101:22:chipyard.TestHarness.RocketConfig.fir@89177.6]
  assign _T_1 = |meta_clients; // @[MSHR.scala 102:29:chipyard.TestHarness.RocketConfig.fir@89179.8]
  assign _T_2 = ~_T_1; // @[MSHR.scala 102:15:chipyard.TestHarness.RocketConfig.fir@89180.8]
  assign _T_4 = _T_2 | reset; // @[MSHR.scala 102:14:chipyard.TestHarness.RocketConfig.fir@89182.8]
  assign _T_5 = ~_T_4; // @[MSHR.scala 102:14:chipyard.TestHarness.RocketConfig.fir@89183.8]
  assign _T_6 = ~meta_dirty; // @[MSHR.scala 103:15:chipyard.TestHarness.RocketConfig.fir@89188.8]
  assign _T_8 = _T_6 | reset; // @[MSHR.scala 103:14:chipyard.TestHarness.RocketConfig.fir@89190.8]
  assign _T_9 = ~_T_8; // @[MSHR.scala 103:14:chipyard.TestHarness.RocketConfig.fir@89191.8]
  assign _T_10 = meta_state == 2'h1; // @[MSHR.scala 105:22:chipyard.TestHarness.RocketConfig.fir@89197.6]
  assign _T_15 = meta_state == 2'h2; // @[MSHR.scala 108:22:chipyard.TestHarness.RocketConfig.fir@89208.6]
  assign _T_18 = _T_1 | reset; // @[MSHR.scala 109:14:chipyard.TestHarness.RocketConfig.fir@89212.8]
  assign _T_19 = ~_T_18; // @[MSHR.scala 109:14:chipyard.TestHarness.RocketConfig.fir@89213.8]
  assign _T_21 = meta_clients - 1'h1; // @[MSHR.scala 110:45:chipyard.TestHarness.RocketConfig.fir@89219.8]
  assign _T_22 = meta_clients & _T_21; // @[MSHR.scala 110:29:chipyard.TestHarness.RocketConfig.fir@89220.8]
  assign _T_23 = ~_T_22; // @[MSHR.scala 110:57:chipyard.TestHarness.RocketConfig.fir@89221.8]
  assign _T_25 = _T_23 | reset; // @[MSHR.scala 110:14:chipyard.TestHarness.RocketConfig.fir@89223.8]
  assign _T_26 = ~_T_25; // @[MSHR.scala 110:14:chipyard.TestHarness.RocketConfig.fir@89224.8]
  assign _T_27 = meta_state == 2'h3; // @[MSHR.scala 112:22:chipyard.TestHarness.RocketConfig.fir@89230.6]
  assign _T_28 = meta_state != 2'h0; // @[MSHR.scala 152:34:chipyard.TestHarness.RocketConfig.fir@89259.4]
  assign _T_29 = meta_valid & _T_28; // @[MSHR.scala 152:20:chipyard.TestHarness.RocketConfig.fir@89260.4]
  assign _T_30 = io_nestedwb_set == request_set; // @[MSHR.scala 153:25:chipyard.TestHarness.RocketConfig.fir@89261.4]
  assign _T_31 = _T_29 & _T_30; // @[MSHR.scala 152:46:chipyard.TestHarness.RocketConfig.fir@89262.4]
  assign _T_32 = io_nestedwb_tag == meta_tag; // @[MSHR.scala 153:60:chipyard.TestHarness.RocketConfig.fir@89263.4]
  assign _T_33 = _T_31 & _T_32; // @[MSHR.scala 153:41:chipyard.TestHarness.RocketConfig.fir@89264.4]
  assign _GEN_0 = io_nestedwb_b_clr_dirty ? 1'h0 : meta_dirty; // @[MSHR.scala 154:36:chipyard.TestHarness.RocketConfig.fir@89266.6]
  assign _GEN_1 = io_nestedwb_c_set_dirty | _GEN_0; // @[MSHR.scala 155:36:chipyard.TestHarness.RocketConfig.fir@89269.6]
  assign _GEN_4 = _T_33 ? _GEN_1 : meta_dirty; // @[MSHR.scala 153:74:chipyard.TestHarness.RocketConfig.fir@89265.4]
  assign _T_34 = ~meta_valid; // @[MSHR.scala 165:28:chipyard.TestHarness.RocketConfig.fir@89283.4]
  assign _T_35 = ~w_releaseack; // @[MSHR.scala 165:45:chipyard.TestHarness.RocketConfig.fir@89284.4]
  assign _T_36 = ~w_rprobeacklast; // @[MSHR.scala 165:62:chipyard.TestHarness.RocketConfig.fir@89285.4]
  assign _T_37 = _T_35 | _T_36; // @[MSHR.scala 165:59:chipyard.TestHarness.RocketConfig.fir@89286.4]
  assign _T_38 = ~w_pprobeacklast; // @[MSHR.scala 165:82:chipyard.TestHarness.RocketConfig.fir@89287.4]
  assign _T_39 = _T_37 | _T_38; // @[MSHR.scala 165:79:chipyard.TestHarness.RocketConfig.fir@89288.4]
  assign _T_40 = ~w_grantfirst; // @[MSHR.scala 165:103:chipyard.TestHarness.RocketConfig.fir@89289.4]
  assign _T_41 = _T_39 & _T_40; // @[MSHR.scala 165:100:chipyard.TestHarness.RocketConfig.fir@89290.4]
  assign _T_43 = meta_valid & w_releaseack; // @[MSHR.scala 166:39:chipyard.TestHarness.RocketConfig.fir@89293.4]
  assign _T_44 = _T_43 & w_rprobeacklast; // @[MSHR.scala 166:55:chipyard.TestHarness.RocketConfig.fir@89294.4]
  assign _T_45 = _T_44 & w_pprobeacklast; // @[MSHR.scala 166:74:chipyard.TestHarness.RocketConfig.fir@89295.4]
  assign _T_49 = ~w_rprobeackfirst; // @[MSHR.scala 170:43:chipyard.TestHarness.RocketConfig.fir@89301.4]
  assign _T_50 = ~w_pprobeackfirst; // @[MSHR.scala 170:64:chipyard.TestHarness.RocketConfig.fir@89302.4]
  assign _T_51 = _T_49 | _T_50; // @[MSHR.scala 170:61:chipyard.TestHarness.RocketConfig.fir@89303.4]
  assign _T_53 = _T_51 | _T_40; // @[MSHR.scala 170:82:chipyard.TestHarness.RocketConfig.fir@89305.4]
  assign _T_55 = ~io_status_bits_nestB; // @[MSHR.scala 176:11:chipyard.TestHarness.RocketConfig.fir@89308.4]
  assign _T_56 = ~io_status_bits_blockB; // @[MSHR.scala 176:36:chipyard.TestHarness.RocketConfig.fir@89309.4]
  assign _T_57 = _T_55 | _T_56; // @[MSHR.scala 176:33:chipyard.TestHarness.RocketConfig.fir@89310.4]
  assign _T_59 = _T_57 | reset; // @[MSHR.scala 176:10:chipyard.TestHarness.RocketConfig.fir@89312.4]
  assign _T_60 = ~_T_59; // @[MSHR.scala 176:10:chipyard.TestHarness.RocketConfig.fir@89313.4]
  assign _T_61 = ~io_status_bits_nestC; // @[MSHR.scala 177:11:chipyard.TestHarness.RocketConfig.fir@89318.4]
  assign _T_62 = ~io_status_bits_blockC; // @[MSHR.scala 177:36:chipyard.TestHarness.RocketConfig.fir@89319.4]
  assign _T_63 = _T_61 | _T_62; // @[MSHR.scala 177:33:chipyard.TestHarness.RocketConfig.fir@89320.4]
  assign _T_65 = _T_63 | reset; // @[MSHR.scala 177:10:chipyard.TestHarness.RocketConfig.fir@89322.4]
  assign _T_66 = ~_T_65; // @[MSHR.scala 177:10:chipyard.TestHarness.RocketConfig.fir@89323.4]
  assign _T_67 = w_rprobeacklast & w_releaseack; // @[MSHR.scala 180:33:chipyard.TestHarness.RocketConfig.fir@89328.4]
  assign _T_68 = _T_67 & w_grantlast; // @[MSHR.scala 180:49:chipyard.TestHarness.RocketConfig.fir@89329.4]
  assign _T_69 = _T_68 & w_pprobeacklast; // @[MSHR.scala 180:64:chipyard.TestHarness.RocketConfig.fir@89330.4]
  assign no_wait = _T_69 & w_grantack; // @[MSHR.scala 180:83:chipyard.TestHarness.RocketConfig.fir@89331.4]
  assign _T_70 = ~s_acquire; // @[MSHR.scala 181:31:chipyard.TestHarness.RocketConfig.fir@89332.4]
  assign _T_71 = _T_70 & s_release; // @[MSHR.scala 181:42:chipyard.TestHarness.RocketConfig.fir@89333.4]
  assign _T_73 = ~s_rprobe; // @[MSHR.scala 182:31:chipyard.TestHarness.RocketConfig.fir@89336.4]
  assign _T_74 = ~s_pprobe; // @[MSHR.scala 182:44:chipyard.TestHarness.RocketConfig.fir@89337.4]
  assign _T_76 = ~s_release; // @[MSHR.scala 183:32:chipyard.TestHarness.RocketConfig.fir@89340.4]
  assign _T_77 = _T_76 & w_rprobeackfirst; // @[MSHR.scala 183:43:chipyard.TestHarness.RocketConfig.fir@89341.4]
  assign _T_81 = ~s_execute; // @[MSHR.scala 184:31:chipyard.TestHarness.RocketConfig.fir@89346.4]
  assign _T_82 = _T_81 & w_pprobeack; // @[MSHR.scala 184:42:chipyard.TestHarness.RocketConfig.fir@89347.4]
  assign _T_84 = ~s_grantack; // @[MSHR.scala 185:31:chipyard.TestHarness.RocketConfig.fir@89350.4]
  assign _T_86 = ~s_flush; // @[MSHR.scala 186:31:chipyard.TestHarness.RocketConfig.fir@89353.4]
  assign _T_90 = ~s_writeback; // @[MSHR.scala 187:70:chipyard.TestHarness.RocketConfig.fir@89358.4]
  assign _T_91 = _T_90 & no_wait; // @[MSHR.scala 187:83:chipyard.TestHarness.RocketConfig.fir@89359.4]
  assign _T_93 = io_schedule_bits_a_valid | io_schedule_bits_b_valid; // @[MSHR.scala 189:49:chipyard.TestHarness.RocketConfig.fir@89363.4]
  assign _T_94 = _T_93 | io_schedule_bits_c_valid; // @[MSHR.scala 189:77:chipyard.TestHarness.RocketConfig.fir@89364.4]
  assign _T_95 = _T_94 | io_schedule_bits_d_valid; // @[MSHR.scala 189:105:chipyard.TestHarness.RocketConfig.fir@89365.4]
  assign _T_96 = _T_95 | io_schedule_bits_e_valid; // @[MSHR.scala 190:49:chipyard.TestHarness.RocketConfig.fir@89366.4]
  assign _T_97 = _T_96 | io_schedule_bits_x_valid; // @[MSHR.scala 190:77:chipyard.TestHarness.RocketConfig.fir@89367.4]
  assign _GEN_7 = w_rprobeackfirst | s_release; // @[MSHR.scala 196:35:chipyard.TestHarness.RocketConfig.fir@89372.6]
  assign _T_99 = s_release & s_pprobe; // @[MSHR.scala 198:21:chipyard.TestHarness.RocketConfig.fir@89376.6]
  assign _GEN_8 = _T_99 | s_acquire; // @[MSHR.scala 198:35:chipyard.TestHarness.RocketConfig.fir@89377.6]
  assign _GEN_9 = w_releaseack | s_flush; // @[MSHR.scala 199:35:chipyard.TestHarness.RocketConfig.fir@89380.6]
  assign _GEN_11 = w_grantfirst | s_grantack; // @[MSHR.scala 201:35:chipyard.TestHarness.RocketConfig.fir@89386.6]
  assign _T_100 = w_pprobeack & w_grant; // @[MSHR.scala 202:23:chipyard.TestHarness.RocketConfig.fir@89389.6]
  assign _GEN_12 = _T_100 | s_execute; // @[MSHR.scala 202:35:chipyard.TestHarness.RocketConfig.fir@89390.6]
  assign _GEN_13 = no_wait | s_writeback; // @[MSHR.scala 203:35:chipyard.TestHarness.RocketConfig.fir@89393.6]
  assign _GEN_14 = no_wait ? 1'h0 : request_valid; // @[MSHR.scala 205:20:chipyard.TestHarness.RocketConfig.fir@89396.6]
  assign _GEN_15 = no_wait ? 1'h0 : meta_valid; // @[MSHR.scala 205:20:chipyard.TestHarness.RocketConfig.fir@89396.6]
  assign _GEN_16 = io_schedule_ready | s_rprobe; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  assign _GEN_17 = io_schedule_ready ? _GEN_7 : s_release; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  assign _GEN_18 = io_schedule_ready | s_pprobe; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  assign _GEN_19 = io_schedule_ready ? _GEN_8 : s_acquire; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  assign _GEN_20 = io_schedule_ready ? _GEN_9 : s_flush; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  assign _GEN_22 = io_schedule_ready ? _GEN_11 : s_grantack; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  assign _GEN_23 = io_schedule_ready ? _GEN_12 : s_execute; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  assign _GEN_24 = io_schedule_ready ? _GEN_13 : s_writeback; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  assign _GEN_25 = io_schedule_ready ? _GEN_14 : request_valid; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  assign _GEN_26 = io_schedule_ready ? _GEN_15 : meta_valid; // @[MSHR.scala 194:28:chipyard.TestHarness.RocketConfig.fir@89370.4]
  assign req_clientBit = request_source == 3'h0; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@89404.4]
  assign _T_102 = ~request_opcode[2]; // @[Parameters.scala 265:5:chipyard.TestHarness.RocketConfig.fir@89406.4]
  assign _T_103 = request_opcode == 3'h5; // @[Parameters.scala 266:13:chipyard.TestHarness.RocketConfig.fir@89407.4]
  assign _T_104 = request_param == 3'h1; // @[Parameters.scala 266:42:chipyard.TestHarness.RocketConfig.fir@89408.4]
  assign _T_105 = _T_103 & _T_104; // @[Parameters.scala 266:33:chipyard.TestHarness.RocketConfig.fir@89409.4]
  assign _T_106 = _T_102 | _T_105; // @[Parameters.scala 265:16:chipyard.TestHarness.RocketConfig.fir@89410.4]
  assign _T_107 = request_opcode == 3'h6; // @[Parameters.scala 267:14:chipyard.TestHarness.RocketConfig.fir@89411.4]
  assign _T_108 = request_opcode == 3'h7; // @[Parameters.scala 267:52:chipyard.TestHarness.RocketConfig.fir@89412.4]
  assign _T_109 = _T_107 | _T_108; // @[Parameters.scala 267:42:chipyard.TestHarness.RocketConfig.fir@89413.4]
  assign _T_110 = request_param != 3'h0; // @[Parameters.scala 267:89:chipyard.TestHarness.RocketConfig.fir@89414.4]
  assign _T_111 = _T_109 & _T_110; // @[Parameters.scala 267:80:chipyard.TestHarness.RocketConfig.fir@89415.4]
  assign req_needT = _T_106 | _T_111; // @[Parameters.scala 266:70:chipyard.TestHarness.RocketConfig.fir@89416.4]
  assign _T_116 = _T_2 & _T_27; // @[MSHR.scala 218:67:chipyard.TestHarness.RocketConfig.fir@89423.4]
  assign _T_117 = meta_hit ? _T_116 : gotT; // @[MSHR.scala 218:40:chipyard.TestHarness.RocketConfig.fir@89424.4]
  assign req_promoteT = _T_109 & _T_117; // @[MSHR.scala 218:34:chipyard.TestHarness.RocketConfig.fir@89425.4]
  assign _T_120 = meta_dirty | request_opcode[0]; // @[MSHR.scala 221:48:chipyard.TestHarness.RocketConfig.fir@89429.6]
  assign _T_121 = request_param != 3'h3; // @[MSHR.scala 222:55:chipyard.TestHarness.RocketConfig.fir@89431.6]
  assign _T_123 = _T_121 & _T_15; // @[MSHR.scala 222:64:chipyard.TestHarness.RocketConfig.fir@89433.6]
  assign _T_124 = _T_123 ? 2'h3 : meta_state; // @[MSHR.scala 222:40:chipyard.TestHarness.RocketConfig.fir@89434.6]
  assign _T_126 = request_param == 3'h2; // @[Parameters.scala 278:43:chipyard.TestHarness.RocketConfig.fir@89437.6]
  assign _T_127 = _T_104 | _T_126; // @[Parameters.scala 278:34:chipyard.TestHarness.RocketConfig.fir@89438.6]
  assign _T_128 = request_param == 3'h5; // @[Parameters.scala 278:75:chipyard.TestHarness.RocketConfig.fir@89439.6]
  assign _T_129 = _T_127 | _T_128; // @[Parameters.scala 278:66:chipyard.TestHarness.RocketConfig.fir@89440.6]
  assign _T_130 = _T_129 & req_clientBit; // @[MSHR.scala 223:56:chipyard.TestHarness.RocketConfig.fir@89441.6]
  assign _T_131 = ~_T_130; // @[MSHR.scala 223:52:chipyard.TestHarness.RocketConfig.fir@89442.6]
  assign _T_132 = meta_clients & _T_131; // @[MSHR.scala 223:50:chipyard.TestHarness.RocketConfig.fir@89443.6]
  assign _T_134 = ~probes_toN; // @[MSHR.scala 229:54:chipyard.TestHarness.RocketConfig.fir@89453.10]
  assign _T_135 = meta_clients & _T_134; // @[MSHR.scala 229:52:chipyard.TestHarness.RocketConfig.fir@89454.10]
  assign _GEN_27 = meta_hit ? 1'h0 : meta_dirty; // @[MSHR.scala 226:21:chipyard.TestHarness.RocketConfig.fir@89450.8]
  assign _GEN_28 = meta_hit ? 2'h0 : meta_state; // @[MSHR.scala 226:21:chipyard.TestHarness.RocketConfig.fir@89450.8]
  assign _GEN_29 = meta_hit ? _T_135 : meta_clients; // @[MSHR.scala 226:21:chipyard.TestHarness.RocketConfig.fir@89450.8]
  assign _T_136 = meta_hit & meta_dirty; // @[MSHR.scala 233:45:chipyard.TestHarness.RocketConfig.fir@89460.8]
  assign _T_139 = _T_136 | _T_102; // @[MSHR.scala 233:60:chipyard.TestHarness.RocketConfig.fir@89463.8]
  assign _T_140 = _T_109 ? 2'h2 : 2'h3; // @[MSHR.scala 235:40:chipyard.TestHarness.RocketConfig.fir@89465.8]
  assign _T_141 = ~meta_hit; // @[MSHR.scala 236:41:chipyard.TestHarness.RocketConfig.fir@89466.8]
  assign _T_143 = gotT ? _T_140 : 2'h1; // @[MSHR.scala 236:55:chipyard.TestHarness.RocketConfig.fir@89468.8]
  assign _T_144 = _T_2 & _T_109; // @[MSHR.scala 241:72:chipyard.TestHarness.RocketConfig.fir@89469.8]
  assign _T_145 = _T_144 ? 2'h2 : 2'h3; // @[MSHR.scala 241:55:chipyard.TestHarness.RocketConfig.fir@89470.8]
  assign _T_146 = 2'h1 == meta_state; // @[Mux.scala 80:60:chipyard.TestHarness.RocketConfig.fir@89471.8]
  assign _T_148 = 2'h2 == meta_state; // @[Mux.scala 80:60:chipyard.TestHarness.RocketConfig.fir@89473.8]
  assign _T_149 = _T_148 ? 2'h3 : 2'h1; // @[Mux.scala 80:57:chipyard.TestHarness.RocketConfig.fir@89474.8]
  assign _T_150 = 2'h3 == meta_state; // @[Mux.scala 80:60:chipyard.TestHarness.RocketConfig.fir@89475.8]
  assign _T_151 = _T_150 ? _T_145 : _T_149; // @[Mux.scala 80:57:chipyard.TestHarness.RocketConfig.fir@89476.8]
  assign _T_152 = _T_141 ? _T_143 : _T_151; // @[MSHR.scala 236:40:chipyard.TestHarness.RocketConfig.fir@89477.8]
  assign _T_153 = req_needT ? _T_140 : _T_152; // @[MSHR.scala 234:38:chipyard.TestHarness.RocketConfig.fir@89478.8]
  assign _T_156 = meta_hit & _T_135; // @[MSHR.scala 242:40:chipyard.TestHarness.RocketConfig.fir@89482.8]
  assign _T_157 = _T_109 & req_clientBit; // @[MSHR.scala 243:40:chipyard.TestHarness.RocketConfig.fir@89483.8]
  assign _T_158 = _T_156 | _T_157; // @[MSHR.scala 242:88:chipyard.TestHarness.RocketConfig.fir@89484.8]
  assign _GEN_30 = request_control ? _GEN_27 : _T_139; // @[MSHR.scala 225:57:chipyard.TestHarness.RocketConfig.fir@89449.6]
  assign _GEN_31 = request_control ? _GEN_28 : _T_153; // @[MSHR.scala 225:57:chipyard.TestHarness.RocketConfig.fir@89449.6]
  assign _GEN_32 = request_control ? _GEN_29 : _T_158; // @[MSHR.scala 225:57:chipyard.TestHarness.RocketConfig.fir@89449.6]
  assign _GEN_33 = request_control ? 1'h0 : 1'h1; // @[MSHR.scala 225:57:chipyard.TestHarness.RocketConfig.fir@89449.6]
  assign _GEN_34 = request_control ? meta_tag : request_tag; // @[MSHR.scala 225:57:chipyard.TestHarness.RocketConfig.fir@89449.6]
  assign _GEN_35 = request_prio_2 ? _T_120 : _GEN_30; // @[MSHR.scala 220:54:chipyard.TestHarness.RocketConfig.fir@89427.4]
  assign _GEN_36 = request_prio_2 ? _T_124 : _GEN_31; // @[MSHR.scala 220:54:chipyard.TestHarness.RocketConfig.fir@89427.4]
  assign _GEN_37 = request_prio_2 ? _T_132 : _GEN_32; // @[MSHR.scala 220:54:chipyard.TestHarness.RocketConfig.fir@89427.4]
  assign _GEN_38 = request_prio_2 | _GEN_33; // @[MSHR.scala 220:54:chipyard.TestHarness.RocketConfig.fir@89427.4]
  assign final_meta_writeback_tag = request_prio_2 ? meta_tag : _GEN_34; // @[MSHR.scala 220:54:chipyard.TestHarness.RocketConfig.fir@89427.4]
  assign _T_161 = _T_34 | _T_10; // @[MSHR.scala 251:27:chipyard.TestHarness.RocketConfig.fir@89493.8]
  assign _T_163 = _T_161 | reset; // @[MSHR.scala 251:14:chipyard.TestHarness.RocketConfig.fir@89495.8]
  assign _T_164 = ~_T_163; // @[MSHR.scala 251:14:chipyard.TestHarness.RocketConfig.fir@89496.8]
  assign _GEN_42 = meta_hit ? 2'h1 : 2'h0; // @[MSHR.scala 249:21:chipyard.TestHarness.RocketConfig.fir@89490.6]
  assign final_meta_writeback_hit = bad_grant ? meta_hit : _GEN_38; // @[MSHR.scala 248:20:chipyard.TestHarness.RocketConfig.fir@89489.4]
  assign final_meta_writeback_dirty = bad_grant ? 1'h0 : _GEN_35; // @[MSHR.scala 248:20:chipyard.TestHarness.RocketConfig.fir@89489.4]
  assign final_meta_writeback_state = bad_grant ? _GEN_42 : _GEN_36; // @[MSHR.scala 248:20:chipyard.TestHarness.RocketConfig.fir@89489.4]
  assign final_meta_writeback_clients = bad_grant ? _T_156 : _GEN_37; // @[MSHR.scala 248:20:chipyard.TestHarness.RocketConfig.fir@89489.4]
  assign _T_167 = meta_clients & req_clientBit; // @[MSHR.scala 273:47:chipyard.TestHarness.RocketConfig.fir@89521.4]
  assign _T_168 = |_T_167; // @[MSHR.scala 273:64:chipyard.TestHarness.RocketConfig.fir@89522.4]
  assign honour_BtoT = meta_hit & _T_168; // @[MSHR.scala 273:30:chipyard.TestHarness.RocketConfig.fir@89523.4]
  assign _T_169 = meta_hit & request_prio_0; // @[MSHR.scala 276:38:chipyard.TestHarness.RocketConfig.fir@89524.4]
  assign _T_173 = request_opcode == 3'h4; // @[Parameters.scala 275:87:chipyard.TestHarness.RocketConfig.fir@89528.4]
  assign _T_174 = _T_109 | _T_173; // @[Parameters.scala 275:77:chipyard.TestHarness.RocketConfig.fir@89529.4]
  assign _T_175 = _T_169 & _T_174; // @[MSHR.scala 276:57:chipyard.TestHarness.RocketConfig.fir@89530.4]
  assign excluded_client = _T_175 & req_clientBit; // @[MSHR.scala 276:28:chipyard.TestHarness.RocketConfig.fir@89531.4]
  assign _T_176 = meta_hit ? 2'h2 : 2'h1; // @[MSHR.scala 279:56:chipyard.TestHarness.RocketConfig.fir@89534.4]
  assign _T_177 = req_needT ? _T_176 : 2'h0; // @[MSHR.scala 279:41:chipyard.TestHarness.RocketConfig.fir@89535.4]
  assign _T_178 = request_size != 3'h6; // @[MSHR.scala 280:51:chipyard.TestHarness.RocketConfig.fir@89537.4]
  assign _T_179 = request_opcode == 3'h0; // @[MSHR.scala 281:55:chipyard.TestHarness.RocketConfig.fir@89538.4]
  assign _T_181 = _T_179 | _T_108; // @[MSHR.scala 281:71:chipyard.TestHarness.RocketConfig.fir@89540.4]
  assign _T_182 = ~_T_181; // @[MSHR.scala 281:38:chipyard.TestHarness.RocketConfig.fir@89541.4]
  assign _T_185 = req_needT ? 2'h2 : 2'h1; // @[MSHR.scala 283:97:chipyard.TestHarness.RocketConfig.fir@89546.4]
  assign _T_186 = request_prio_1 ? request_param : {{1'd0}, _T_185}; // @[MSHR.scala 283:61:chipyard.TestHarness.RocketConfig.fir@89547.4]
  assign _T_190 = ~excluded_client; // @[MSHR.scala 286:53:chipyard.TestHarness.RocketConfig.fir@89554.4]
  assign _T_191 = meta_clients & _T_190; // @[MSHR.scala 286:51:chipyard.TestHarness.RocketConfig.fir@89555.4]
  assign _T_195 = ~_T_109; // @[MSHR.scala 295:42:chipyard.TestHarness.RocketConfig.fir@89568.4]
  assign _T_197 = req_promoteT ? 2'h1 : 2'h0; // @[MSHR.scala 297:53:chipyard.TestHarness.RocketConfig.fir@89571.4]
  assign _T_198 = honour_BtoT ? 2'h2 : 2'h1; // @[MSHR.scala 298:53:chipyard.TestHarness.RocketConfig.fir@89572.4]
  assign _T_199 = 3'h0 == request_param; // @[Mux.scala 80:60:chipyard.TestHarness.RocketConfig.fir@89573.4]
  assign _T_200 = _T_199 ? {{1'd0}, _T_197} : 3'h0; // @[Mux.scala 80:57:chipyard.TestHarness.RocketConfig.fir@89574.4]
  assign _T_201 = 3'h2 == request_param; // @[Mux.scala 80:60:chipyard.TestHarness.RocketConfig.fir@89575.4]
  assign _T_202 = _T_201 ? {{1'd0}, _T_198} : _T_200; // @[Mux.scala 80:57:chipyard.TestHarness.RocketConfig.fir@89576.4]
  assign _T_203 = 3'h1 == request_param; // @[Mux.scala 80:60:chipyard.TestHarness.RocketConfig.fir@89577.4]
  assign _T_204 = _T_203 ? 3'h1 : _T_202; // @[Mux.scala 80:57:chipyard.TestHarness.RocketConfig.fir@89578.4]
  assign _T_212 = _T_1 ? 1'h0 : 1'h1; // @[MSHR.scala 315:32:chipyard.TestHarness.RocketConfig.fir@89600.6]
  assign _T_214 = meta_dirty ? 2'h2 : 2'h3; // @[MSHR.scala 316:32:chipyard.TestHarness.RocketConfig.fir@89606.8]
  assign _T_216 = meta_dirty ? 3'h4 : 3'h5; // @[MSHR.scala 317:39:chipyard.TestHarness.RocketConfig.fir@89612.10]
  assign _T_217 = meta_dirty ? 3'h6 : 3'h7; // @[MSHR.scala 317:76:chipyard.TestHarness.RocketConfig.fir@89613.10]
  assign _T_218 = _T_1 ? _T_216 : _T_217; // @[MSHR.scala 317:32:chipyard.TestHarness.RocketConfig.fir@89614.10]
  assign _GEN_49 = _T_150 ? {{1'd0}, _T_218} : 4'h8; // @[Conditional.scala 39:67:chipyard.TestHarness.RocketConfig.fir@89611.8]
  assign _GEN_50 = _T_148 ? {{2'd0}, _T_214} : _GEN_49; // @[Conditional.scala 39:67:chipyard.TestHarness.RocketConfig.fir@89605.6]
  assign _GEN_51 = _T_146 ? {{3'd0}, _T_212} : _GEN_50; // @[Conditional.scala 40:58:chipyard.TestHarness.RocketConfig.fir@89599.4]
  assign _T_220 = ~_T_141; // @[MSHR.scala 320:11:chipyard.TestHarness.RocketConfig.fir@89622.4]
  assign evict = _T_220 ? 4'h8 : _GEN_51; // @[MSHR.scala 320:17:chipyard.TestHarness.RocketConfig.fir@89623.4]
  assign before_ = _T_141 ? 4'h8 : _GEN_51; // @[MSHR.scala 320:17:chipyard.TestHarness.RocketConfig.fir@89654.4]
  assign _T_232 = |final_meta_writeback_clients; // @[MSHR.scala 312:27:chipyard.TestHarness.RocketConfig.fir@89659.4]
  assign _T_233 = 2'h1 == final_meta_writeback_state; // @[Conditional.scala 37:30:chipyard.TestHarness.RocketConfig.fir@89660.4]
  assign _T_234 = _T_232 ? 1'h0 : 1'h1; // @[MSHR.scala 315:32:chipyard.TestHarness.RocketConfig.fir@89662.6]
  assign _T_235 = 2'h2 == final_meta_writeback_state; // @[Conditional.scala 37:30:chipyard.TestHarness.RocketConfig.fir@89666.6]
  assign _T_236 = final_meta_writeback_dirty ? 2'h2 : 2'h3; // @[MSHR.scala 316:32:chipyard.TestHarness.RocketConfig.fir@89668.8]
  assign _T_237 = 2'h3 == final_meta_writeback_state; // @[Conditional.scala 37:30:chipyard.TestHarness.RocketConfig.fir@89672.8]
  assign _T_238 = final_meta_writeback_dirty ? 3'h4 : 3'h5; // @[MSHR.scala 317:39:chipyard.TestHarness.RocketConfig.fir@89674.10]
  assign _T_239 = final_meta_writeback_dirty ? 3'h6 : 3'h7; // @[MSHR.scala 317:76:chipyard.TestHarness.RocketConfig.fir@89675.10]
  assign _T_240 = _T_232 ? _T_238 : _T_239; // @[MSHR.scala 317:32:chipyard.TestHarness.RocketConfig.fir@89676.10]
  assign _GEN_59 = _T_237 ? {{1'd0}, _T_240} : 4'h8; // @[Conditional.scala 39:67:chipyard.TestHarness.RocketConfig.fir@89673.8]
  assign _GEN_60 = _T_235 ? {{2'd0}, _T_236} : _GEN_59; // @[Conditional.scala 39:67:chipyard.TestHarness.RocketConfig.fir@89667.6]
  assign after = _T_233 ? {{3'd0}, _T_234} : _GEN_60; // @[Conditional.scala 40:58:chipyard.TestHarness.RocketConfig.fir@89661.4]
  assign _T_245 = _T_77 & io_schedule_ready; // @[MSHR.scala 360:42:chipyard.TestHarness.RocketConfig.fir@89690.4]
  assign _T_246 = evict == 4'h1; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89692.6]
  assign _T_247 = ~_T_246; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89693.6]
  assign _T_249 = _T_247 | reset; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89695.6]
  assign _T_250 = ~_T_249; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89696.6]
  assign _T_251 = before_ == 4'h1; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89701.6]
  assign _T_252 = ~_T_251; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89702.6]
  assign _T_254 = _T_252 | reset; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89704.6]
  assign _T_255 = ~_T_254; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89705.6]
  assign _T_256 = evict == 4'h0; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89710.6]
  assign _T_257 = ~_T_256; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89711.6]
  assign _T_259 = _T_257 | reset; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89713.6]
  assign _T_260 = ~_T_259; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89714.6]
  assign _T_261 = before_ == 4'h0; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89719.6]
  assign _T_262 = ~_T_261; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89720.6]
  assign _T_264 = _T_262 | reset; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89722.6]
  assign _T_265 = ~_T_264; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89723.6]
  assign _T_267 = before_ == 4'h7; // @[MSHR.scala 363:13:chipyard.TestHarness.RocketConfig.fir@89729.6]
  assign _T_269 = before_ == 4'h5; // @[MSHR.scala 364:13:chipyard.TestHarness.RocketConfig.fir@89731.6]
  assign _T_271 = before_ == 4'h4; // @[MSHR.scala 365:13:chipyard.TestHarness.RocketConfig.fir@89733.6]
  assign _T_273 = before_ == 4'h6; // @[MSHR.scala 366:13:chipyard.TestHarness.RocketConfig.fir@89735.6]
  assign _T_275 = before_ == 4'h3; // @[MSHR.scala 367:13:chipyard.TestHarness.RocketConfig.fir@89737.6]
  assign _T_277 = before_ == 4'h2; // @[MSHR.scala 368:13:chipyard.TestHarness.RocketConfig.fir@89739.6]
  assign _T_280 = _T_91 & io_schedule_ready; // @[MSHR.scala 371:35:chipyard.TestHarness.RocketConfig.fir@89743.4]
  assign _T_281 = before_ == 4'h8; // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89745.6]
  assign _T_282 = after == 4'h1; // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89746.6]
  assign _T_283 = _T_281 & _T_282; // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89747.6]
  assign _T_284 = ~_T_283; // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89748.6]
  assign _T_286 = _T_284 | reset; // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89750.6]
  assign _T_287 = ~_T_286; // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89751.6]
  assign _T_289 = after == 4'h0; // @[MSHR.scala 373:15:chipyard.TestHarness.RocketConfig.fir@89757.6]
  assign _T_290 = _T_281 & _T_289; // @[MSHR.scala 373:15:chipyard.TestHarness.RocketConfig.fir@89758.6]
  assign _T_291 = ~_T_290; // @[MSHR.scala 373:15:chipyard.TestHarness.RocketConfig.fir@89759.6]
  assign _T_293 = _T_291 | reset; // @[MSHR.scala 373:15:chipyard.TestHarness.RocketConfig.fir@89761.6]
  assign _T_294 = ~_T_293; // @[MSHR.scala 373:15:chipyard.TestHarness.RocketConfig.fir@89762.6]
  assign _T_296 = after == 4'h7; // @[MSHR.scala 374:15:chipyard.TestHarness.RocketConfig.fir@89768.6]
  assign _T_299 = after == 4'h5; // @[MSHR.scala 375:15:chipyard.TestHarness.RocketConfig.fir@89771.6]
  assign _T_300 = _T_281 & _T_299; // @[MSHR.scala 375:15:chipyard.TestHarness.RocketConfig.fir@89772.6]
  assign _T_301 = ~_T_300; // @[MSHR.scala 375:15:chipyard.TestHarness.RocketConfig.fir@89773.6]
  assign _T_303 = _T_301 | reset; // @[MSHR.scala 375:15:chipyard.TestHarness.RocketConfig.fir@89775.6]
  assign _T_304 = ~_T_303; // @[MSHR.scala 375:15:chipyard.TestHarness.RocketConfig.fir@89776.6]
  assign _T_306 = after == 4'h4; // @[MSHR.scala 376:15:chipyard.TestHarness.RocketConfig.fir@89782.6]
  assign _T_307 = _T_281 & _T_306; // @[MSHR.scala 376:15:chipyard.TestHarness.RocketConfig.fir@89783.6]
  assign _T_308 = ~_T_307; // @[MSHR.scala 376:15:chipyard.TestHarness.RocketConfig.fir@89784.6]
  assign _T_310 = _T_308 | reset; // @[MSHR.scala 376:15:chipyard.TestHarness.RocketConfig.fir@89786.6]
  assign _T_311 = ~_T_310; // @[MSHR.scala 376:15:chipyard.TestHarness.RocketConfig.fir@89787.6]
  assign _T_313 = after == 4'h6; // @[MSHR.scala 377:15:chipyard.TestHarness.RocketConfig.fir@89793.6]
  assign _T_316 = after == 4'h3; // @[MSHR.scala 378:15:chipyard.TestHarness.RocketConfig.fir@89796.6]
  assign _T_319 = after == 4'h2; // @[MSHR.scala 379:15:chipyard.TestHarness.RocketConfig.fir@89799.6]
  assign _T_320 = _T_281 & _T_319; // @[MSHR.scala 379:15:chipyard.TestHarness.RocketConfig.fir@89800.6]
  assign _T_321 = ~_T_320; // @[MSHR.scala 379:15:chipyard.TestHarness.RocketConfig.fir@89801.6]
  assign _T_323 = _T_321 | reset; // @[MSHR.scala 379:15:chipyard.TestHarness.RocketConfig.fir@89803.6]
  assign _T_324 = ~_T_323; // @[MSHR.scala 379:15:chipyard.TestHarness.RocketConfig.fir@89804.6]
  assign _T_326 = after == 4'h8; // @[MSHR.scala 381:15:chipyard.TestHarness.RocketConfig.fir@89810.6]
  assign _T_327 = _T_251 & _T_326; // @[MSHR.scala 381:15:chipyard.TestHarness.RocketConfig.fir@89811.6]
  assign _T_328 = ~_T_327; // @[MSHR.scala 381:15:chipyard.TestHarness.RocketConfig.fir@89812.6]
  assign _T_330 = _T_328 | reset; // @[MSHR.scala 381:15:chipyard.TestHarness.RocketConfig.fir@89814.6]
  assign _T_331 = ~_T_330; // @[MSHR.scala 381:15:chipyard.TestHarness.RocketConfig.fir@89815.6]
  assign _T_334 = _T_251 & _T_289; // @[MSHR.scala 382:15:chipyard.TestHarness.RocketConfig.fir@89822.6]
  assign _T_335 = ~_T_334; // @[MSHR.scala 382:15:chipyard.TestHarness.RocketConfig.fir@89823.6]
  assign _T_337 = _T_335 | reset; // @[MSHR.scala 382:15:chipyard.TestHarness.RocketConfig.fir@89825.6]
  assign _T_338 = ~_T_337; // @[MSHR.scala 382:15:chipyard.TestHarness.RocketConfig.fir@89826.6]
  assign _T_341 = _T_251 & _T_296; // @[MSHR.scala 383:15:chipyard.TestHarness.RocketConfig.fir@89833.6]
  assign _T_342 = ~_T_341; // @[MSHR.scala 383:15:chipyard.TestHarness.RocketConfig.fir@89834.6]
  assign _T_344 = _T_342 | reset; // @[MSHR.scala 383:15:chipyard.TestHarness.RocketConfig.fir@89836.6]
  assign _T_345 = ~_T_344; // @[MSHR.scala 383:15:chipyard.TestHarness.RocketConfig.fir@89837.6]
  assign _T_348 = _T_251 & _T_299; // @[MSHR.scala 384:15:chipyard.TestHarness.RocketConfig.fir@89844.6]
  assign _T_349 = ~_T_348; // @[MSHR.scala 384:15:chipyard.TestHarness.RocketConfig.fir@89845.6]
  assign _T_351 = _T_349 | reset; // @[MSHR.scala 384:15:chipyard.TestHarness.RocketConfig.fir@89847.6]
  assign _T_352 = ~_T_351; // @[MSHR.scala 384:15:chipyard.TestHarness.RocketConfig.fir@89848.6]
  assign _T_355 = _T_251 & _T_306; // @[MSHR.scala 385:15:chipyard.TestHarness.RocketConfig.fir@89855.6]
  assign _T_356 = ~_T_355; // @[MSHR.scala 385:15:chipyard.TestHarness.RocketConfig.fir@89856.6]
  assign _T_358 = _T_356 | reset; // @[MSHR.scala 385:15:chipyard.TestHarness.RocketConfig.fir@89858.6]
  assign _T_359 = ~_T_358; // @[MSHR.scala 385:15:chipyard.TestHarness.RocketConfig.fir@89859.6]
  assign _T_362 = _T_251 & _T_313; // @[MSHR.scala 386:15:chipyard.TestHarness.RocketConfig.fir@89866.6]
  assign _T_363 = ~_T_362; // @[MSHR.scala 386:15:chipyard.TestHarness.RocketConfig.fir@89867.6]
  assign _T_365 = _T_363 | reset; // @[MSHR.scala 386:15:chipyard.TestHarness.RocketConfig.fir@89869.6]
  assign _T_366 = ~_T_365; // @[MSHR.scala 386:15:chipyard.TestHarness.RocketConfig.fir@89870.6]
  assign _T_369 = _T_251 & _T_316; // @[MSHR.scala 387:15:chipyard.TestHarness.RocketConfig.fir@89877.6]
  assign _T_370 = ~_T_369; // @[MSHR.scala 387:15:chipyard.TestHarness.RocketConfig.fir@89878.6]
  assign _T_372 = _T_370 | reset; // @[MSHR.scala 387:15:chipyard.TestHarness.RocketConfig.fir@89880.6]
  assign _T_373 = ~_T_372; // @[MSHR.scala 387:15:chipyard.TestHarness.RocketConfig.fir@89881.6]
  assign _T_376 = _T_251 & _T_319; // @[MSHR.scala 388:15:chipyard.TestHarness.RocketConfig.fir@89888.6]
  assign _T_377 = ~_T_376; // @[MSHR.scala 388:15:chipyard.TestHarness.RocketConfig.fir@89889.6]
  assign _T_379 = _T_377 | reset; // @[MSHR.scala 388:15:chipyard.TestHarness.RocketConfig.fir@89891.6]
  assign _T_380 = ~_T_379; // @[MSHR.scala 388:15:chipyard.TestHarness.RocketConfig.fir@89892.6]
  assign _T_383 = _T_261 & _T_326; // @[MSHR.scala 390:15:chipyard.TestHarness.RocketConfig.fir@89899.6]
  assign _T_384 = ~_T_383; // @[MSHR.scala 390:15:chipyard.TestHarness.RocketConfig.fir@89900.6]
  assign _T_386 = _T_384 | reset; // @[MSHR.scala 390:15:chipyard.TestHarness.RocketConfig.fir@89902.6]
  assign _T_387 = ~_T_386; // @[MSHR.scala 390:15:chipyard.TestHarness.RocketConfig.fir@89903.6]
  assign _T_390 = _T_261 & _T_282; // @[MSHR.scala 391:15:chipyard.TestHarness.RocketConfig.fir@89910.6]
  assign _T_391 = ~_T_390; // @[MSHR.scala 391:15:chipyard.TestHarness.RocketConfig.fir@89911.6]
  assign _T_393 = _T_391 | reset; // @[MSHR.scala 391:15:chipyard.TestHarness.RocketConfig.fir@89913.6]
  assign _T_394 = ~_T_393; // @[MSHR.scala 391:15:chipyard.TestHarness.RocketConfig.fir@89914.6]
  assign _T_397 = _T_261 & _T_296; // @[MSHR.scala 392:15:chipyard.TestHarness.RocketConfig.fir@89921.6]
  assign _T_398 = ~_T_397; // @[MSHR.scala 392:15:chipyard.TestHarness.RocketConfig.fir@89922.6]
  assign _T_400 = _T_398 | reset; // @[MSHR.scala 392:15:chipyard.TestHarness.RocketConfig.fir@89924.6]
  assign _T_401 = ~_T_400; // @[MSHR.scala 392:15:chipyard.TestHarness.RocketConfig.fir@89925.6]
  assign _T_404 = _T_261 & _T_299; // @[MSHR.scala 393:15:chipyard.TestHarness.RocketConfig.fir@89932.6]
  assign _T_405 = ~_T_404; // @[MSHR.scala 393:15:chipyard.TestHarness.RocketConfig.fir@89933.6]
  assign _T_407 = _T_405 | reset; // @[MSHR.scala 393:15:chipyard.TestHarness.RocketConfig.fir@89935.6]
  assign _T_408 = ~_T_407; // @[MSHR.scala 393:15:chipyard.TestHarness.RocketConfig.fir@89936.6]
  assign _T_411 = _T_261 & _T_313; // @[MSHR.scala 394:15:chipyard.TestHarness.RocketConfig.fir@89943.6]
  assign _T_412 = ~_T_411; // @[MSHR.scala 394:15:chipyard.TestHarness.RocketConfig.fir@89944.6]
  assign _T_414 = _T_412 | reset; // @[MSHR.scala 394:15:chipyard.TestHarness.RocketConfig.fir@89946.6]
  assign _T_415 = ~_T_414; // @[MSHR.scala 394:15:chipyard.TestHarness.RocketConfig.fir@89947.6]
  assign _T_418 = _T_261 & _T_306; // @[MSHR.scala 395:15:chipyard.TestHarness.RocketConfig.fir@89954.6]
  assign _T_419 = ~_T_418; // @[MSHR.scala 395:15:chipyard.TestHarness.RocketConfig.fir@89955.6]
  assign _T_421 = _T_419 | reset; // @[MSHR.scala 395:15:chipyard.TestHarness.RocketConfig.fir@89957.6]
  assign _T_422 = ~_T_421; // @[MSHR.scala 395:15:chipyard.TestHarness.RocketConfig.fir@89958.6]
  assign _T_425 = _T_261 & _T_316; // @[MSHR.scala 396:15:chipyard.TestHarness.RocketConfig.fir@89965.6]
  assign _T_426 = ~_T_425; // @[MSHR.scala 396:15:chipyard.TestHarness.RocketConfig.fir@89966.6]
  assign _T_428 = _T_426 | reset; // @[MSHR.scala 396:15:chipyard.TestHarness.RocketConfig.fir@89968.6]
  assign _T_429 = ~_T_428; // @[MSHR.scala 396:15:chipyard.TestHarness.RocketConfig.fir@89969.6]
  assign _T_432 = _T_261 & _T_319; // @[MSHR.scala 397:15:chipyard.TestHarness.RocketConfig.fir@89976.6]
  assign _T_433 = ~_T_432; // @[MSHR.scala 397:15:chipyard.TestHarness.RocketConfig.fir@89977.6]
  assign _T_435 = _T_433 | reset; // @[MSHR.scala 397:15:chipyard.TestHarness.RocketConfig.fir@89979.6]
  assign _T_436 = ~_T_435; // @[MSHR.scala 397:15:chipyard.TestHarness.RocketConfig.fir@89980.6]
  assign _T_439 = _T_267 & _T_326; // @[MSHR.scala 399:15:chipyard.TestHarness.RocketConfig.fir@89987.6]
  assign _T_440 = ~_T_439; // @[MSHR.scala 399:15:chipyard.TestHarness.RocketConfig.fir@89988.6]
  assign _T_442 = _T_440 | reset; // @[MSHR.scala 399:15:chipyard.TestHarness.RocketConfig.fir@89990.6]
  assign _T_443 = ~_T_442; // @[MSHR.scala 399:15:chipyard.TestHarness.RocketConfig.fir@89991.6]
  assign _T_446 = _T_267 & _T_282; // @[MSHR.scala 400:15:chipyard.TestHarness.RocketConfig.fir@89998.6]
  assign _T_447 = ~_T_446; // @[MSHR.scala 400:15:chipyard.TestHarness.RocketConfig.fir@89999.6]
  assign _T_449 = _T_447 | reset; // @[MSHR.scala 400:15:chipyard.TestHarness.RocketConfig.fir@90001.6]
  assign _T_450 = ~_T_449; // @[MSHR.scala 400:15:chipyard.TestHarness.RocketConfig.fir@90002.6]
  assign _T_453 = _T_267 & _T_289; // @[MSHR.scala 401:15:chipyard.TestHarness.RocketConfig.fir@90009.6]
  assign _T_454 = ~_T_453; // @[MSHR.scala 401:15:chipyard.TestHarness.RocketConfig.fir@90010.6]
  assign _T_456 = _T_454 | reset; // @[MSHR.scala 401:15:chipyard.TestHarness.RocketConfig.fir@90012.6]
  assign _T_457 = ~_T_456; // @[MSHR.scala 401:15:chipyard.TestHarness.RocketConfig.fir@90013.6]
  assign _T_460 = _T_267 & _T_299; // @[MSHR.scala 402:15:chipyard.TestHarness.RocketConfig.fir@90020.6]
  assign _T_461 = ~_T_460; // @[MSHR.scala 402:15:chipyard.TestHarness.RocketConfig.fir@90021.6]
  assign _T_463 = _T_461 | reset; // @[MSHR.scala 402:15:chipyard.TestHarness.RocketConfig.fir@90023.6]
  assign _T_464 = ~_T_463; // @[MSHR.scala 402:15:chipyard.TestHarness.RocketConfig.fir@90024.6]
  assign _T_470 = _T_267 & _T_306; // @[MSHR.scala 404:15:chipyard.TestHarness.RocketConfig.fir@90034.6]
  assign _T_471 = ~_T_470; // @[MSHR.scala 404:15:chipyard.TestHarness.RocketConfig.fir@90035.6]
  assign _T_473 = _T_471 | reset; // @[MSHR.scala 404:15:chipyard.TestHarness.RocketConfig.fir@90037.6]
  assign _T_474 = ~_T_473; // @[MSHR.scala 404:15:chipyard.TestHarness.RocketConfig.fir@90038.6]
  assign _T_480 = _T_267 & _T_319; // @[MSHR.scala 406:15:chipyard.TestHarness.RocketConfig.fir@90048.6]
  assign _T_481 = ~_T_480; // @[MSHR.scala 406:15:chipyard.TestHarness.RocketConfig.fir@90049.6]
  assign _T_483 = _T_481 | reset; // @[MSHR.scala 406:15:chipyard.TestHarness.RocketConfig.fir@90051.6]
  assign _T_484 = ~_T_483; // @[MSHR.scala 406:15:chipyard.TestHarness.RocketConfig.fir@90052.6]
  assign _T_487 = _T_269 & _T_326; // @[MSHR.scala 408:15:chipyard.TestHarness.RocketConfig.fir@90059.6]
  assign _T_488 = ~_T_487; // @[MSHR.scala 408:15:chipyard.TestHarness.RocketConfig.fir@90060.6]
  assign _T_490 = _T_488 | reset; // @[MSHR.scala 408:15:chipyard.TestHarness.RocketConfig.fir@90062.6]
  assign _T_491 = ~_T_490; // @[MSHR.scala 408:15:chipyard.TestHarness.RocketConfig.fir@90063.6]
  assign _T_494 = _T_269 & _T_282; // @[MSHR.scala 409:15:chipyard.TestHarness.RocketConfig.fir@90070.6]
  assign _T_495 = ~_T_494; // @[MSHR.scala 409:15:chipyard.TestHarness.RocketConfig.fir@90071.6]
  assign _T_497 = _T_495 | reset; // @[MSHR.scala 409:15:chipyard.TestHarness.RocketConfig.fir@90073.6]
  assign _T_498 = ~_T_497; // @[MSHR.scala 409:15:chipyard.TestHarness.RocketConfig.fir@90074.6]
  assign _T_501 = _T_269 & _T_289; // @[MSHR.scala 410:15:chipyard.TestHarness.RocketConfig.fir@90081.6]
  assign _T_502 = ~_T_501; // @[MSHR.scala 410:15:chipyard.TestHarness.RocketConfig.fir@90082.6]
  assign _T_504 = _T_502 | reset; // @[MSHR.scala 410:15:chipyard.TestHarness.RocketConfig.fir@90084.6]
  assign _T_505 = ~_T_504; // @[MSHR.scala 410:15:chipyard.TestHarness.RocketConfig.fir@90085.6]
  assign _T_514 = _T_269 & _T_306; // @[MSHR.scala 413:15:chipyard.TestHarness.RocketConfig.fir@90098.6]
  assign _T_515 = ~_T_514; // @[MSHR.scala 413:15:chipyard.TestHarness.RocketConfig.fir@90099.6]
  assign _T_517 = _T_515 | reset; // @[MSHR.scala 413:15:chipyard.TestHarness.RocketConfig.fir@90101.6]
  assign _T_518 = ~_T_517; // @[MSHR.scala 413:15:chipyard.TestHarness.RocketConfig.fir@90102.6]
  assign _T_524 = _T_269 & _T_319; // @[MSHR.scala 415:15:chipyard.TestHarness.RocketConfig.fir@90112.6]
  assign _T_525 = ~_T_524; // @[MSHR.scala 415:15:chipyard.TestHarness.RocketConfig.fir@90113.6]
  assign _T_527 = _T_525 | reset; // @[MSHR.scala 415:15:chipyard.TestHarness.RocketConfig.fir@90115.6]
  assign _T_528 = ~_T_527; // @[MSHR.scala 415:15:chipyard.TestHarness.RocketConfig.fir@90116.6]
  assign _T_531 = _T_273 & _T_326; // @[MSHR.scala 417:15:chipyard.TestHarness.RocketConfig.fir@90123.6]
  assign _T_532 = ~_T_531; // @[MSHR.scala 417:15:chipyard.TestHarness.RocketConfig.fir@90124.6]
  assign _T_534 = _T_532 | reset; // @[MSHR.scala 417:15:chipyard.TestHarness.RocketConfig.fir@90126.6]
  assign _T_535 = ~_T_534; // @[MSHR.scala 417:15:chipyard.TestHarness.RocketConfig.fir@90127.6]
  assign _T_538 = _T_273 & _T_282; // @[MSHR.scala 418:15:chipyard.TestHarness.RocketConfig.fir@90134.6]
  assign _T_539 = ~_T_538; // @[MSHR.scala 418:15:chipyard.TestHarness.RocketConfig.fir@90135.6]
  assign _T_541 = _T_539 | reset; // @[MSHR.scala 418:15:chipyard.TestHarness.RocketConfig.fir@90137.6]
  assign _T_542 = ~_T_541; // @[MSHR.scala 418:15:chipyard.TestHarness.RocketConfig.fir@90138.6]
  assign _T_545 = _T_273 & _T_289; // @[MSHR.scala 419:15:chipyard.TestHarness.RocketConfig.fir@90145.6]
  assign _T_546 = ~_T_545; // @[MSHR.scala 419:15:chipyard.TestHarness.RocketConfig.fir@90146.6]
  assign _T_548 = _T_546 | reset; // @[MSHR.scala 419:15:chipyard.TestHarness.RocketConfig.fir@90148.6]
  assign _T_549 = ~_T_548; // @[MSHR.scala 419:15:chipyard.TestHarness.RocketConfig.fir@90149.6]
  assign _T_552 = _T_273 & _T_296; // @[MSHR.scala 420:15:chipyard.TestHarness.RocketConfig.fir@90156.6]
  assign _T_553 = ~_T_552; // @[MSHR.scala 420:15:chipyard.TestHarness.RocketConfig.fir@90157.6]
  assign _T_555 = _T_553 | reset; // @[MSHR.scala 420:15:chipyard.TestHarness.RocketConfig.fir@90159.6]
  assign _T_556 = ~_T_555; // @[MSHR.scala 420:15:chipyard.TestHarness.RocketConfig.fir@90160.6]
  assign _T_559 = _T_273 & _T_299; // @[MSHR.scala 421:15:chipyard.TestHarness.RocketConfig.fir@90167.6]
  assign _T_560 = ~_T_559; // @[MSHR.scala 421:15:chipyard.TestHarness.RocketConfig.fir@90168.6]
  assign _T_562 = _T_560 | reset; // @[MSHR.scala 421:15:chipyard.TestHarness.RocketConfig.fir@90170.6]
  assign _T_563 = ~_T_562; // @[MSHR.scala 421:15:chipyard.TestHarness.RocketConfig.fir@90171.6]
  assign _T_566 = _T_273 & _T_306; // @[MSHR.scala 422:15:chipyard.TestHarness.RocketConfig.fir@90178.6]
  assign _T_567 = ~_T_566; // @[MSHR.scala 422:15:chipyard.TestHarness.RocketConfig.fir@90179.6]
  assign _T_569 = _T_567 | reset; // @[MSHR.scala 422:15:chipyard.TestHarness.RocketConfig.fir@90181.6]
  assign _T_570 = ~_T_569; // @[MSHR.scala 422:15:chipyard.TestHarness.RocketConfig.fir@90182.6]
  assign _T_573 = _T_273 & _T_316; // @[MSHR.scala 423:15:chipyard.TestHarness.RocketConfig.fir@90189.6]
  assign _T_574 = ~_T_573; // @[MSHR.scala 423:15:chipyard.TestHarness.RocketConfig.fir@90190.6]
  assign _T_576 = _T_574 | reset; // @[MSHR.scala 423:15:chipyard.TestHarness.RocketConfig.fir@90192.6]
  assign _T_577 = ~_T_576; // @[MSHR.scala 423:15:chipyard.TestHarness.RocketConfig.fir@90193.6]
  assign _T_583 = _T_271 & _T_326; // @[MSHR.scala 426:15:chipyard.TestHarness.RocketConfig.fir@90203.6]
  assign _T_584 = ~_T_583; // @[MSHR.scala 426:15:chipyard.TestHarness.RocketConfig.fir@90204.6]
  assign _T_586 = _T_584 | reset; // @[MSHR.scala 426:15:chipyard.TestHarness.RocketConfig.fir@90206.6]
  assign _T_587 = ~_T_586; // @[MSHR.scala 426:15:chipyard.TestHarness.RocketConfig.fir@90207.6]
  assign _T_590 = _T_271 & _T_282; // @[MSHR.scala 427:15:chipyard.TestHarness.RocketConfig.fir@90214.6]
  assign _T_591 = ~_T_590; // @[MSHR.scala 427:15:chipyard.TestHarness.RocketConfig.fir@90215.6]
  assign _T_593 = _T_591 | reset; // @[MSHR.scala 427:15:chipyard.TestHarness.RocketConfig.fir@90217.6]
  assign _T_594 = ~_T_593; // @[MSHR.scala 427:15:chipyard.TestHarness.RocketConfig.fir@90218.6]
  assign _T_597 = _T_271 & _T_289; // @[MSHR.scala 428:15:chipyard.TestHarness.RocketConfig.fir@90225.6]
  assign _T_598 = ~_T_597; // @[MSHR.scala 428:15:chipyard.TestHarness.RocketConfig.fir@90226.6]
  assign _T_600 = _T_598 | reset; // @[MSHR.scala 428:15:chipyard.TestHarness.RocketConfig.fir@90228.6]
  assign _T_601 = ~_T_600; // @[MSHR.scala 428:15:chipyard.TestHarness.RocketConfig.fir@90229.6]
  assign _T_604 = _T_271 & _T_296; // @[MSHR.scala 429:15:chipyard.TestHarness.RocketConfig.fir@90236.6]
  assign _T_605 = ~_T_604; // @[MSHR.scala 429:15:chipyard.TestHarness.RocketConfig.fir@90237.6]
  assign _T_607 = _T_605 | reset; // @[MSHR.scala 429:15:chipyard.TestHarness.RocketConfig.fir@90239.6]
  assign _T_608 = ~_T_607; // @[MSHR.scala 429:15:chipyard.TestHarness.RocketConfig.fir@90240.6]
  assign _T_611 = _T_271 & _T_299; // @[MSHR.scala 430:15:chipyard.TestHarness.RocketConfig.fir@90247.6]
  assign _T_612 = ~_T_611; // @[MSHR.scala 430:15:chipyard.TestHarness.RocketConfig.fir@90248.6]
  assign _T_614 = _T_612 | reset; // @[MSHR.scala 430:15:chipyard.TestHarness.RocketConfig.fir@90250.6]
  assign _T_615 = ~_T_614; // @[MSHR.scala 430:15:chipyard.TestHarness.RocketConfig.fir@90251.6]
  assign _T_621 = _T_271 & _T_316; // @[MSHR.scala 432:15:chipyard.TestHarness.RocketConfig.fir@90261.6]
  assign _T_622 = ~_T_621; // @[MSHR.scala 432:15:chipyard.TestHarness.RocketConfig.fir@90262.6]
  assign _T_624 = _T_622 | reset; // @[MSHR.scala 432:15:chipyard.TestHarness.RocketConfig.fir@90264.6]
  assign _T_625 = ~_T_624; // @[MSHR.scala 432:15:chipyard.TestHarness.RocketConfig.fir@90265.6]
  assign _T_631 = _T_275 & _T_326; // @[MSHR.scala 435:15:chipyard.TestHarness.RocketConfig.fir@90275.6]
  assign _T_632 = ~_T_631; // @[MSHR.scala 435:15:chipyard.TestHarness.RocketConfig.fir@90276.6]
  assign _T_634 = _T_632 | reset; // @[MSHR.scala 435:15:chipyard.TestHarness.RocketConfig.fir@90278.6]
  assign _T_635 = ~_T_634; // @[MSHR.scala 435:15:chipyard.TestHarness.RocketConfig.fir@90279.6]
  assign _T_638 = _T_275 & _T_282; // @[MSHR.scala 436:15:chipyard.TestHarness.RocketConfig.fir@90286.6]
  assign _T_639 = ~_T_638; // @[MSHR.scala 436:15:chipyard.TestHarness.RocketConfig.fir@90287.6]
  assign _T_641 = _T_639 | reset; // @[MSHR.scala 436:15:chipyard.TestHarness.RocketConfig.fir@90289.6]
  assign _T_642 = ~_T_641; // @[MSHR.scala 436:15:chipyard.TestHarness.RocketConfig.fir@90290.6]
  assign _T_645 = _T_275 & _T_289; // @[MSHR.scala 437:15:chipyard.TestHarness.RocketConfig.fir@90297.6]
  assign _T_646 = ~_T_645; // @[MSHR.scala 437:15:chipyard.TestHarness.RocketConfig.fir@90298.6]
  assign _T_648 = _T_646 | reset; // @[MSHR.scala 437:15:chipyard.TestHarness.RocketConfig.fir@90300.6]
  assign _T_649 = ~_T_648; // @[MSHR.scala 437:15:chipyard.TestHarness.RocketConfig.fir@90301.6]
  assign _T_667 = _T_277 & _T_326; // @[MSHR.scala 444:15:chipyard.TestHarness.RocketConfig.fir@90323.6]
  assign _T_668 = ~_T_667; // @[MSHR.scala 444:15:chipyard.TestHarness.RocketConfig.fir@90324.6]
  assign _T_670 = _T_668 | reset; // @[MSHR.scala 444:15:chipyard.TestHarness.RocketConfig.fir@90326.6]
  assign _T_671 = ~_T_670; // @[MSHR.scala 444:15:chipyard.TestHarness.RocketConfig.fir@90327.6]
  assign _T_674 = _T_277 & _T_282; // @[MSHR.scala 445:15:chipyard.TestHarness.RocketConfig.fir@90334.6]
  assign _T_675 = ~_T_674; // @[MSHR.scala 445:15:chipyard.TestHarness.RocketConfig.fir@90335.6]
  assign _T_677 = _T_675 | reset; // @[MSHR.scala 445:15:chipyard.TestHarness.RocketConfig.fir@90337.6]
  assign _T_678 = ~_T_677; // @[MSHR.scala 445:15:chipyard.TestHarness.RocketConfig.fir@90338.6]
  assign _T_681 = _T_277 & _T_289; // @[MSHR.scala 446:15:chipyard.TestHarness.RocketConfig.fir@90345.6]
  assign _T_682 = ~_T_681; // @[MSHR.scala 446:15:chipyard.TestHarness.RocketConfig.fir@90346.6]
  assign _T_684 = _T_682 | reset; // @[MSHR.scala 446:15:chipyard.TestHarness.RocketConfig.fir@90348.6]
  assign _T_685 = ~_T_684; // @[MSHR.scala 446:15:chipyard.TestHarness.RocketConfig.fir@90349.6]
  assign _T_688 = _T_277 & _T_296; // @[MSHR.scala 447:15:chipyard.TestHarness.RocketConfig.fir@90356.6]
  assign _T_689 = ~_T_688; // @[MSHR.scala 447:15:chipyard.TestHarness.RocketConfig.fir@90357.6]
  assign _T_691 = _T_689 | reset; // @[MSHR.scala 447:15:chipyard.TestHarness.RocketConfig.fir@90359.6]
  assign _T_692 = ~_T_691; // @[MSHR.scala 447:15:chipyard.TestHarness.RocketConfig.fir@90360.6]
  assign _T_695 = _T_277 & _T_299; // @[MSHR.scala 448:15:chipyard.TestHarness.RocketConfig.fir@90367.6]
  assign _T_696 = ~_T_695; // @[MSHR.scala 448:15:chipyard.TestHarness.RocketConfig.fir@90368.6]
  assign _T_698 = _T_696 | reset; // @[MSHR.scala 448:15:chipyard.TestHarness.RocketConfig.fir@90370.6]
  assign _T_699 = ~_T_698; // @[MSHR.scala 448:15:chipyard.TestHarness.RocketConfig.fir@90371.6]
  assign _T_708 = _T_277 & _T_316; // @[MSHR.scala 451:15:chipyard.TestHarness.RocketConfig.fir@90384.6]
  assign _T_709 = ~_T_708; // @[MSHR.scala 451:15:chipyard.TestHarness.RocketConfig.fir@90385.6]
  assign _T_711 = _T_709 | reset; // @[MSHR.scala 451:15:chipyard.TestHarness.RocketConfig.fir@90387.6]
  assign _T_712 = ~_T_711; // @[MSHR.scala 451:15:chipyard.TestHarness.RocketConfig.fir@90388.6]
  assign probe_bit = io_sinkc_bits_source == 3'h0; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@90394.4]
  assign _T_713 = probes_done | probe_bit; // @[MSHR.scala 456:33:chipyard.TestHarness.RocketConfig.fir@90395.4]
  assign last_probe = _T_713 == _T_191; // @[MSHR.scala 456:46:chipyard.TestHarness.RocketConfig.fir@90398.4]
  assign _T_716 = io_sinkc_bits_param == 3'h1; // @[Parameters.scala 278:11:chipyard.TestHarness.RocketConfig.fir@90399.4]
  assign _T_717 = io_sinkc_bits_param == 3'h2; // @[Parameters.scala 278:43:chipyard.TestHarness.RocketConfig.fir@90400.4]
  assign _T_718 = _T_716 | _T_717; // @[Parameters.scala 278:34:chipyard.TestHarness.RocketConfig.fir@90401.4]
  assign _T_719 = io_sinkc_bits_param == 3'h5; // @[Parameters.scala 278:75:chipyard.TestHarness.RocketConfig.fir@90402.4]
  assign probe_toN = _T_718 | _T_719; // @[Parameters.scala 278:66:chipyard.TestHarness.RocketConfig.fir@90403.4]
  assign _T_726 = probe_toN & probe_bit; // @[MSHR.scala 465:35:chipyard.TestHarness.RocketConfig.fir@90412.6]
  assign _T_727 = probes_toN | _T_726; // @[MSHR.scala 465:30:chipyard.TestHarness.RocketConfig.fir@90413.6]
  assign _T_730 = w_rprobeackfirst | last_probe; // @[MSHR.scala 467:42:chipyard.TestHarness.RocketConfig.fir@90418.6]
  assign _T_731 = last_probe & io_sinkc_bits_last; // @[MSHR.scala 468:55:chipyard.TestHarness.RocketConfig.fir@90420.6]
  assign _T_732 = w_rprobeacklast | _T_731; // @[MSHR.scala 468:40:chipyard.TestHarness.RocketConfig.fir@90421.6]
  assign _T_733 = w_pprobeackfirst | last_probe; // @[MSHR.scala 469:42:chipyard.TestHarness.RocketConfig.fir@90423.6]
  assign _T_735 = w_pprobeacklast | _T_731; // @[MSHR.scala 470:40:chipyard.TestHarness.RocketConfig.fir@90426.6]
  assign _T_736 = request_offset == 6'h0; // @[MSHR.scala 472:77:chipyard.TestHarness.RocketConfig.fir@90428.6]
  assign _T_737 = io_sinkc_bits_last | _T_736; // @[MSHR.scala 472:59:chipyard.TestHarness.RocketConfig.fir@90429.6]
  assign _T_738 = last_probe & _T_737; // @[MSHR.scala 472:36:chipyard.TestHarness.RocketConfig.fir@90430.6]
  assign _T_739 = w_pprobeack | _T_738; // @[MSHR.scala 473:32:chipyard.TestHarness.RocketConfig.fir@90431.6]
  assign _T_744 = io_sinkc_bits_tag == meta_tag; // @[MSHR.scala 477:55:chipyard.TestHarness.RocketConfig.fir@90437.6]
  assign _T_745 = _T_28 & _T_744; // @[MSHR.scala 477:34:chipyard.TestHarness.RocketConfig.fir@90438.6]
  assign _T_746 = _T_745 & io_sinkc_bits_data; // @[MSHR.scala 477:68:chipyard.TestHarness.RocketConfig.fir@90439.6]
  assign _GEN_63 = _T_746 | _GEN_4; // @[MSHR.scala 477:91:chipyard.TestHarness.RocketConfig.fir@90440.6]
  assign _GEN_67 = io_sinkc_valid ? _T_730 : w_rprobeackfirst; // @[MSHR.scala 458:49:chipyard.TestHarness.RocketConfig.fir@90404.4]
  assign _GEN_68 = io_sinkc_valid ? _T_732 : w_rprobeacklast; // @[MSHR.scala 458:49:chipyard.TestHarness.RocketConfig.fir@90404.4]
  assign _GEN_69 = io_sinkc_valid ? _T_733 : w_pprobeackfirst; // @[MSHR.scala 458:49:chipyard.TestHarness.RocketConfig.fir@90404.4]
  assign _GEN_70 = io_sinkc_valid ? _T_735 : w_pprobeacklast; // @[MSHR.scala 458:49:chipyard.TestHarness.RocketConfig.fir@90404.4]
  assign _GEN_71 = io_sinkc_valid ? _T_739 : w_pprobeack; // @[MSHR.scala 458:49:chipyard.TestHarness.RocketConfig.fir@90404.4]
  assign _T_747 = io_sinkd_bits_opcode == 3'h4; // @[MSHR.scala 480:32:chipyard.TestHarness.RocketConfig.fir@90445.6]
  assign _T_748 = io_sinkd_bits_opcode == 3'h5; // @[MSHR.scala 480:66:chipyard.TestHarness.RocketConfig.fir@90446.6]
  assign _T_749 = _T_747 | _T_748; // @[MSHR.scala 480:42:chipyard.TestHarness.RocketConfig.fir@90447.6]
  assign _T_751 = _T_736 | io_sinkd_bits_last; // @[MSHR.scala 487:45:chipyard.TestHarness.RocketConfig.fir@90454.8]
  assign _T_758 = io_sinkd_bits_param == 3'h0; // @[MSHR.scala 490:35:chipyard.TestHarness.RocketConfig.fir@90462.8]
  assign _T_759 = io_sinkd_bits_opcode == 3'h6; // @[MSHR.scala 492:37:chipyard.TestHarness.RocketConfig.fir@90466.8]
  assign _GEN_73 = _T_759 | w_releaseack; // @[MSHR.scala 492:53:chipyard.TestHarness.RocketConfig.fir@90467.8]
  assign _GEN_75 = _T_749 | w_grantfirst; // @[MSHR.scala 480:81:chipyard.TestHarness.RocketConfig.fir@90448.6]
  assign _GEN_76 = _T_749 ? io_sinkd_bits_last : w_grantlast; // @[MSHR.scala 480:81:chipyard.TestHarness.RocketConfig.fir@90448.6]
  assign _GEN_78 = _T_749 ? _T_751 : w_grant; // @[MSHR.scala 480:81:chipyard.TestHarness.RocketConfig.fir@90448.6]
  assign _GEN_80 = _T_749 ? w_releaseack : _GEN_73; // @[MSHR.scala 480:81:chipyard.TestHarness.RocketConfig.fir@90448.6]
  assign _GEN_82 = io_sinkd_valid ? _GEN_75 : w_grantfirst; // @[MSHR.scala 479:25:chipyard.TestHarness.RocketConfig.fir@90444.4]
  assign _GEN_83 = io_sinkd_valid ? _GEN_76 : w_grantlast; // @[MSHR.scala 479:25:chipyard.TestHarness.RocketConfig.fir@90444.4]
  assign _GEN_85 = io_sinkd_valid ? _GEN_78 : w_grant; // @[MSHR.scala 479:25:chipyard.TestHarness.RocketConfig.fir@90444.4]
  assign _GEN_87 = io_sinkd_valid ? _GEN_80 : w_releaseack; // @[MSHR.scala 479:25:chipyard.TestHarness.RocketConfig.fir@90444.4]
  assign _GEN_88 = io_sinke_valid | w_grantack; // @[MSHR.scala 496:25:chipyard.TestHarness.RocketConfig.fir@90471.4]
  assign _T_760 = io_allocate_valid & io_allocate_bits_repeat; // @[MSHR.scala 502:40:chipyard.TestHarness.RocketConfig.fir@90477.4]
  assign new_meta_dirty = _T_760 ? final_meta_writeback_dirty : io_directory_bits_dirty; // @[MSHR.scala 502:21:chipyard.TestHarness.RocketConfig.fir@90478.4]
  assign new_meta_state = _T_760 ? final_meta_writeback_state : io_directory_bits_state; // @[MSHR.scala 502:21:chipyard.TestHarness.RocketConfig.fir@90478.4]
  assign new_meta_clients = _T_760 ? final_meta_writeback_clients : io_directory_bits_clients; // @[MSHR.scala 502:21:chipyard.TestHarness.RocketConfig.fir@90478.4]
  assign new_meta_hit = _T_760 ? final_meta_writeback_hit : io_directory_bits_hit; // @[MSHR.scala 502:21:chipyard.TestHarness.RocketConfig.fir@90478.4]
  assign new_request_prio_2 = io_allocate_valid ? io_allocate_bits_prio_2 : request_prio_2; // @[MSHR.scala 503:24:chipyard.TestHarness.RocketConfig.fir@90479.4]
  assign new_request_control = io_allocate_valid ? io_allocate_bits_control : request_control; // @[MSHR.scala 503:24:chipyard.TestHarness.RocketConfig.fir@90479.4]
  assign new_request_opcode = io_allocate_valid ? io_allocate_bits_opcode : request_opcode; // @[MSHR.scala 503:24:chipyard.TestHarness.RocketConfig.fir@90479.4]
  assign new_request_param = io_allocate_valid ? io_allocate_bits_param : request_param; // @[MSHR.scala 503:24:chipyard.TestHarness.RocketConfig.fir@90479.4]
  assign new_request_source = io_allocate_valid ? io_allocate_bits_source : request_source; // @[MSHR.scala 503:24:chipyard.TestHarness.RocketConfig.fir@90479.4]
  assign _T_762 = ~new_request_opcode[2]; // @[Parameters.scala 265:5:chipyard.TestHarness.RocketConfig.fir@90481.4]
  assign _T_763 = new_request_opcode == 3'h5; // @[Parameters.scala 266:13:chipyard.TestHarness.RocketConfig.fir@90482.4]
  assign _T_764 = new_request_param == 3'h1; // @[Parameters.scala 266:42:chipyard.TestHarness.RocketConfig.fir@90483.4]
  assign _T_765 = _T_763 & _T_764; // @[Parameters.scala 266:33:chipyard.TestHarness.RocketConfig.fir@90484.4]
  assign _T_766 = _T_762 | _T_765; // @[Parameters.scala 265:16:chipyard.TestHarness.RocketConfig.fir@90485.4]
  assign _T_767 = new_request_opcode == 3'h6; // @[Parameters.scala 267:14:chipyard.TestHarness.RocketConfig.fir@90486.4]
  assign _T_768 = new_request_opcode == 3'h7; // @[Parameters.scala 267:52:chipyard.TestHarness.RocketConfig.fir@90487.4]
  assign _T_769 = _T_767 | _T_768; // @[Parameters.scala 267:42:chipyard.TestHarness.RocketConfig.fir@90488.4]
  assign _T_770 = new_request_param != 3'h0; // @[Parameters.scala 267:89:chipyard.TestHarness.RocketConfig.fir@90489.4]
  assign _T_771 = _T_769 & _T_770; // @[Parameters.scala 267:80:chipyard.TestHarness.RocketConfig.fir@90490.4]
  assign new_needT = _T_766 | _T_771; // @[Parameters.scala 266:70:chipyard.TestHarness.RocketConfig.fir@90491.4]
  assign new_clientBit = new_request_source == 3'h0; // @[Parameters.scala 47:9:chipyard.TestHarness.RocketConfig.fir@90492.4]
  assign _T_775 = new_request_opcode == 3'h4; // @[Parameters.scala 275:87:chipyard.TestHarness.RocketConfig.fir@90496.4]
  assign _T_776 = _T_769 | _T_775; // @[Parameters.scala 275:77:chipyard.TestHarness.RocketConfig.fir@90497.4]
  assign new_skipProbe = _T_776 & new_clientBit; // @[MSHR.scala 506:26:chipyard.TestHarness.RocketConfig.fir@90498.4]
  assign _T_791 = ~_T_282; // @[MSHR.scala 519:11:chipyard.TestHarness.RocketConfig.fir@90534.6]
  assign _T_793 = _T_791 | reset; // @[MSHR.scala 519:11:chipyard.TestHarness.RocketConfig.fir@90536.6]
  assign _T_794 = ~_T_793; // @[MSHR.scala 519:11:chipyard.TestHarness.RocketConfig.fir@90537.6]
  assign _T_796 = ~_T_289; // @[MSHR.scala 520:11:chipyard.TestHarness.RocketConfig.fir@90543.6]
  assign _T_798 = _T_796 | reset; // @[MSHR.scala 520:11:chipyard.TestHarness.RocketConfig.fir@90545.6]
  assign _T_799 = ~_T_798; // @[MSHR.scala 520:11:chipyard.TestHarness.RocketConfig.fir@90546.6]
  assign _T_806 = ~request_valid; // @[MSHR.scala 530:13:chipyard.TestHarness.RocketConfig.fir@90559.6]
  assign _T_807 = io_schedule_ready & io_schedule_valid; // @[Decoupled.scala 40:37:chipyard.TestHarness.RocketConfig.fir@90560.6]
  assign _T_808 = no_wait & _T_807; // @[MSHR.scala 530:40:chipyard.TestHarness.RocketConfig.fir@90561.6]
  assign _T_809 = _T_806 | _T_808; // @[MSHR.scala 530:28:chipyard.TestHarness.RocketConfig.fir@90562.6]
  assign _T_811 = _T_809 | reset; // @[MSHR.scala 530:12:chipyard.TestHarness.RocketConfig.fir@90564.6]
  assign _T_812 = ~_T_811; // @[MSHR.scala 530:12:chipyard.TestHarness.RocketConfig.fir@90565.6]
  assign _GEN_94 = io_allocate_valid | _GEN_25; // @[MSHR.scala 529:28:chipyard.TestHarness.RocketConfig.fir@90558.4]
  assign _T_814 = io_directory_valid | _T_760; // @[MSHR.scala 536:28:chipyard.TestHarness.RocketConfig.fir@90574.4]
  assign _T_817 = ~new_meta_dirty; // @[MSHR.scala 571:38:chipyard.TestHarness.RocketConfig.fir@90606.8]
  assign _T_818 = new_request_opcode[0] & _T_817; // @[MSHR.scala 571:35:chipyard.TestHarness.RocketConfig.fir@90607.8]
  assign _GEN_107 = _T_818 ? 1'h0 : 1'h1; // @[MSHR.scala 571:55:chipyard.TestHarness.RocketConfig.fir@90608.8]
  assign _T_819 = new_request_param == 3'h0; // @[Parameters.scala 281:11:chipyard.TestHarness.RocketConfig.fir@90611.8]
  assign _T_820 = new_request_param == 3'h4; // @[Parameters.scala 281:43:chipyard.TestHarness.RocketConfig.fir@90612.8]
  assign _T_821 = _T_819 | _T_820; // @[Parameters.scala 281:34:chipyard.TestHarness.RocketConfig.fir@90613.8]
  assign _T_822 = new_meta_state == 2'h2; // @[MSHR.scala 575:56:chipyard.TestHarness.RocketConfig.fir@90614.8]
  assign _T_823 = _T_821 & _T_822; // @[MSHR.scala 575:38:chipyard.TestHarness.RocketConfig.fir@90615.8]
  assign _GEN_108 = _T_823 ? 1'h0 : _GEN_107; // @[MSHR.scala 575:67:chipyard.TestHarness.RocketConfig.fir@90616.8]
  assign _T_825 = new_request_param == 3'h2; // @[Parameters.scala 278:43:chipyard.TestHarness.RocketConfig.fir@90620.8]
  assign _T_826 = _T_764 | _T_825; // @[Parameters.scala 278:34:chipyard.TestHarness.RocketConfig.fir@90621.8]
  assign _T_827 = new_request_param == 3'h5; // @[Parameters.scala 278:75:chipyard.TestHarness.RocketConfig.fir@90622.8]
  assign _T_828 = _T_826 | _T_827; // @[Parameters.scala 278:66:chipyard.TestHarness.RocketConfig.fir@90623.8]
  assign _T_829 = new_meta_clients & new_clientBit; // @[MSHR.scala 579:59:chipyard.TestHarness.RocketConfig.fir@90624.8]
  assign _T_831 = _T_828 & _T_829; // @[MSHR.scala 579:38:chipyard.TestHarness.RocketConfig.fir@90626.8]
  assign _GEN_109 = _T_831 ? 1'h0 : _GEN_108; // @[MSHR.scala 579:89:chipyard.TestHarness.RocketConfig.fir@90627.8]
  assign _T_833 = new_meta_hit | reset; // @[MSHR.scala 582:14:chipyard.TestHarness.RocketConfig.fir@90631.8]
  assign _T_834 = ~_T_833; // @[MSHR.scala 582:14:chipyard.TestHarness.RocketConfig.fir@90632.8]
  assign _GEN_110 = new_meta_clients ? 1'h0 : 1'h1; // @[MSHR.scala 592:75:chipyard.TestHarness.RocketConfig.fir@90647.12]
  assign _GEN_111 = new_meta_hit ? 1'h0 : 1'h1; // @[MSHR.scala 588:27:chipyard.TestHarness.RocketConfig.fir@90642.10]
  assign _GEN_112 = new_meta_hit ? _GEN_110 : 1'h1; // @[MSHR.scala 588:27:chipyard.TestHarness.RocketConfig.fir@90642.10]
  assign _T_838 = ~new_meta_hit; // @[MSHR.scala 603:13:chipyard.TestHarness.RocketConfig.fir@90656.10]
  assign _T_839 = new_meta_state != 2'h0; // @[MSHR.scala 603:45:chipyard.TestHarness.RocketConfig.fir@90657.10]
  assign _T_840 = _T_838 & _T_839; // @[MSHR.scala 603:27:chipyard.TestHarness.RocketConfig.fir@90658.10]
  assign _GEN_114 = _T_840 ? 1'h0 : 1'h1; // @[MSHR.scala 603:58:chipyard.TestHarness.RocketConfig.fir@90659.10]
  assign _GEN_115 = _T_840 ? _GEN_110 : 1'h1; // @[MSHR.scala 603:58:chipyard.TestHarness.RocketConfig.fir@90659.10]
  assign _T_844 = new_meta_state == 2'h1; // @[MSHR.scala 614:46:chipyard.TestHarness.RocketConfig.fir@90671.10]
  assign _T_845 = _T_844 & new_needT; // @[MSHR.scala 614:57:chipyard.TestHarness.RocketConfig.fir@90672.10]
  assign _T_846 = _T_838 | _T_845; // @[MSHR.scala 614:27:chipyard.TestHarness.RocketConfig.fir@90673.10]
  assign _GEN_116 = _T_846 ? 1'h0 : 1'h1; // @[MSHR.scala 614:72:chipyard.TestHarness.RocketConfig.fir@90674.10]
  assign _T_848 = new_needT | _T_822; // @[MSHR.scala 624:24:chipyard.TestHarness.RocketConfig.fir@90683.10]
  assign _T_849 = new_meta_hit & _T_848; // @[MSHR.scala 623:55:chipyard.TestHarness.RocketConfig.fir@90684.10]
  assign _T_850 = ~new_skipProbe; // @[MSHR.scala 625:33:chipyard.TestHarness.RocketConfig.fir@90685.10]
  assign _T_851 = new_meta_clients & _T_850; // @[MSHR.scala 625:31:chipyard.TestHarness.RocketConfig.fir@90686.10]
  assign _T_853 = _T_849 & _T_851; // @[MSHR.scala 624:53:chipyard.TestHarness.RocketConfig.fir@90688.10]
  assign _GEN_117 = _T_853 ? 1'h0 : 1'h1; // @[MSHR.scala 625:63:chipyard.TestHarness.RocketConfig.fir@90690.10]
  assign _GEN_118 = _T_853 ? 1'h0 : _GEN_116; // @[MSHR.scala 625:63:chipyard.TestHarness.RocketConfig.fir@90690.10]
  assign _GEN_119 = _T_769 ? 1'h0 : 1'h1; // @[MSHR.scala 633:88:chipyard.TestHarness.RocketConfig.fir@90700.10]
  assign _GEN_120 = _T_769 ? 1'h0 : _GEN_118; // @[MSHR.scala 633:88:chipyard.TestHarness.RocketConfig.fir@90700.10]
  assign _T_860 = _T_762 & new_meta_hit; // @[MSHR.scala 638:36:chipyard.TestHarness.RocketConfig.fir@90706.10]
  assign _T_862 = _T_860 & _T_817; // @[MSHR.scala 638:52:chipyard.TestHarness.RocketConfig.fir@90708.10]
  assign _GEN_121 = _T_862 ? 1'h0 : _GEN_120; // @[MSHR.scala 638:72:chipyard.TestHarness.RocketConfig.fir@90709.10]
  assign _GEN_122 = new_request_control ? 1'h0 : 1'h1; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  assign _GEN_123 = new_request_control ? _GEN_111 : _GEN_114; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  assign _GEN_124 = new_request_control ? _GEN_112 : _GEN_115; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  assign _GEN_126 = new_request_control | _GEN_116; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  assign _GEN_127 = new_request_control | _GEN_121; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  assign _GEN_128 = new_request_control | _GEN_117; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  assign _GEN_129 = new_request_control | _GEN_119; // @[MSHR.scala 585:61:chipyard.TestHarness.RocketConfig.fir@90640.8]
  assign _GEN_130 = new_request_prio_2 ? 1'h0 : new_request_control; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  assign _GEN_131 = new_request_prio_2 ? _GEN_109 : _GEN_127; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  assign _GEN_132 = new_request_prio_2 | _GEN_122; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  assign _GEN_133 = new_request_prio_2 | _GEN_123; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  assign _GEN_134 = new_request_prio_2 | _GEN_124; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  assign _GEN_135 = new_request_prio_2 | _GEN_126; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  assign _GEN_136 = new_request_prio_2 | _GEN_128; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  assign _GEN_137 = new_request_prio_2 | _GEN_129; // @[MSHR.scala 568:60:chipyard.TestHarness.RocketConfig.fir@90603.6]
  assign _GEN_138 = _T_814 | _GEN_26; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_150 = _T_814 ? _GEN_134 : _GEN_16; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_151 = _T_814 ? _GEN_134 : _GEN_67; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_152 = _T_814 ? _GEN_134 : _GEN_68; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_153 = _T_814 ? _GEN_133 : _GEN_17; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_154 = _T_814 ? _GEN_133 : _GEN_87; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_155 = _T_814 ? _GEN_136 : _GEN_18; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_156 = _T_814 ? _GEN_135 : _GEN_19; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_157 = _T_814 ? _GEN_132 : _GEN_20; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_158 = _T_814 ? _GEN_135 : _GEN_82; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_159 = _T_814 ? _GEN_135 : _GEN_83; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_160 = _T_814 ? _GEN_135 : _GEN_85; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_161 = _T_814 ? _GEN_136 : _GEN_69; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_162 = _T_814 ? _GEN_136 : _GEN_70; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_163 = _T_814 ? _GEN_136 : _GEN_71; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_165 = _T_814 ? _GEN_135 : _GEN_22; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_166 = _T_814 ? _GEN_130 : _GEN_23; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_167 = _T_814 ? _GEN_137 : _GEN_88; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign _GEN_168 = _T_814 ? _GEN_131 : _GEN_24; // @[MSHR.scala 536:79:chipyard.TestHarness.RocketConfig.fir@90575.4]
  assign io_status_valid = request_valid; // @[MSHR.scala 161:19:chipyard.TestHarness.RocketConfig.fir@89279.4]
  assign io_status_bits_set = request_set; // @[MSHR.scala 162:25:chipyard.TestHarness.RocketConfig.fir@89280.4]
  assign io_status_bits_tag = request_tag; // @[MSHR.scala 163:25:chipyard.TestHarness.RocketConfig.fir@89281.4]
  assign io_status_bits_way = meta_way; // @[MSHR.scala 164:25:chipyard.TestHarness.RocketConfig.fir@89282.4]
  assign io_status_bits_blockB = _T_34 | _T_41; // @[MSHR.scala 165:25:chipyard.TestHarness.RocketConfig.fir@89292.4]
  assign io_status_bits_nestB = _T_45 & _T_40; // @[MSHR.scala 166:25:chipyard.TestHarness.RocketConfig.fir@89298.4]
  assign io_status_bits_blockC = ~meta_valid; // @[MSHR.scala 169:25:chipyard.TestHarness.RocketConfig.fir@89300.4]
  assign io_status_bits_nestC = meta_valid & _T_53; // @[MSHR.scala 170:25:chipyard.TestHarness.RocketConfig.fir@89307.4]
  assign io_schedule_valid = _T_97 | io_schedule_bits_dir_valid; // @[MSHR.scala 189:21:chipyard.TestHarness.RocketConfig.fir@89369.4]
  assign io_schedule_bits_a_valid = _T_71 & s_pprobe; // @[MSHR.scala 181:28:chipyard.TestHarness.RocketConfig.fir@89335.4]
  assign io_schedule_bits_a_bits_tag = request_tag; // @[MSHR.scala 277:35:chipyard.TestHarness.RocketConfig.fir@89532.4]
  assign io_schedule_bits_a_bits_set = request_set; // @[MSHR.scala 278:35:chipyard.TestHarness.RocketConfig.fir@89533.4]
  assign io_schedule_bits_a_bits_param = {{1'd0}, _T_177}; // @[MSHR.scala 279:35:chipyard.TestHarness.RocketConfig.fir@89536.4]
  assign io_schedule_bits_a_bits_block = _T_178 | _T_182; // @[MSHR.scala 280:35:chipyard.TestHarness.RocketConfig.fir@89543.4]
  assign io_schedule_bits_b_valid = _T_73 | _T_74; // @[MSHR.scala 182:28:chipyard.TestHarness.RocketConfig.fir@89339.4]
  assign io_schedule_bits_b_bits_param = _T_73 ? 3'h2 : _T_186; // @[MSHR.scala 283:35:chipyard.TestHarness.RocketConfig.fir@89549.4]
  assign io_schedule_bits_b_bits_tag = _T_73 ? meta_tag : request_tag; // @[MSHR.scala 284:35:chipyard.TestHarness.RocketConfig.fir@89552.4]
  assign io_schedule_bits_b_bits_set = request_set; // @[MSHR.scala 285:35:chipyard.TestHarness.RocketConfig.fir@89553.4]
  assign io_schedule_bits_b_bits_clients = meta_clients & _T_190; // @[MSHR.scala 286:35:chipyard.TestHarness.RocketConfig.fir@89556.4]
  assign io_schedule_bits_c_valid = _T_76 & w_rprobeackfirst; // @[MSHR.scala 183:28:chipyard.TestHarness.RocketConfig.fir@89345.4]
  assign io_schedule_bits_c_bits_opcode = meta_dirty ? 3'h7 : 3'h6; // @[MSHR.scala 287:35:chipyard.TestHarness.RocketConfig.fir@89558.4]
  assign io_schedule_bits_c_bits_param = _T_10 ? 3'h2 : 3'h1; // @[MSHR.scala 288:35:chipyard.TestHarness.RocketConfig.fir@89561.4]
  assign io_schedule_bits_c_bits_tag = meta_tag; // @[MSHR.scala 290:35:chipyard.TestHarness.RocketConfig.fir@89563.4]
  assign io_schedule_bits_c_bits_set = request_set; // @[MSHR.scala 291:35:chipyard.TestHarness.RocketConfig.fir@89564.4]
  assign io_schedule_bits_c_bits_way = meta_way; // @[MSHR.scala 292:35:chipyard.TestHarness.RocketConfig.fir@89565.4]
  assign io_schedule_bits_c_bits_dirty = meta_dirty; // @[MSHR.scala 293:35:chipyard.TestHarness.RocketConfig.fir@89566.4]
  assign io_schedule_bits_d_valid = _T_82 & w_grant; // @[MSHR.scala 184:28:chipyard.TestHarness.RocketConfig.fir@89349.4]
  assign io_schedule_bits_d_bits_prio_0 = request_prio_0; // @[MSHR.scala 294:35:chipyard.TestHarness.RocketConfig.fir@89567.4]
  assign io_schedule_bits_d_bits_prio_1 = request_prio_1; // @[MSHR.scala 294:35:chipyard.TestHarness.RocketConfig.fir@89567.4]
  assign io_schedule_bits_d_bits_prio_2 = request_prio_2; // @[MSHR.scala 294:35:chipyard.TestHarness.RocketConfig.fir@89567.4]
  assign io_schedule_bits_d_bits_control = request_control; // @[MSHR.scala 294:35:chipyard.TestHarness.RocketConfig.fir@89567.4]
  assign io_schedule_bits_d_bits_opcode = request_opcode; // @[MSHR.scala 294:35:chipyard.TestHarness.RocketConfig.fir@89567.4]
  assign io_schedule_bits_d_bits_param = _T_195 ? request_param : _T_204; // @[MSHR.scala 294:35:chipyard.TestHarness.RocketConfig.fir@89567.4 MSHR.scala 295:35:chipyard.TestHarness.RocketConfig.fir@89580.4]
  assign io_schedule_bits_d_bits_size = request_size; // @[MSHR.scala 294:35:chipyard.TestHarness.RocketConfig.fir@89567.4]
  assign io_schedule_bits_d_bits_source = request_source; // @[MSHR.scala 294:35:chipyard.TestHarness.RocketConfig.fir@89567.4]
  assign io_schedule_bits_d_bits_tag = request_tag; // @[MSHR.scala 294:35:chipyard.TestHarness.RocketConfig.fir@89567.4]
  assign io_schedule_bits_d_bits_offset = request_offset; // @[MSHR.scala 294:35:chipyard.TestHarness.RocketConfig.fir@89567.4]
  assign io_schedule_bits_d_bits_put = request_put; // @[MSHR.scala 294:35:chipyard.TestHarness.RocketConfig.fir@89567.4]
  assign io_schedule_bits_d_bits_set = request_set; // @[MSHR.scala 294:35:chipyard.TestHarness.RocketConfig.fir@89567.4]
  assign io_schedule_bits_d_bits_way = meta_way; // @[MSHR.scala 301:35:chipyard.TestHarness.RocketConfig.fir@89582.4]
  assign io_schedule_bits_d_bits_bad = bad_grant; // @[MSHR.scala 302:35:chipyard.TestHarness.RocketConfig.fir@89583.4]
  assign io_schedule_bits_e_valid = _T_84 & w_grantfirst; // @[MSHR.scala 185:28:chipyard.TestHarness.RocketConfig.fir@89352.4]
  assign io_schedule_bits_e_bits_sink = sink; // @[MSHR.scala 303:35:chipyard.TestHarness.RocketConfig.fir@89584.4]
  assign io_schedule_bits_x_valid = _T_86 & w_releaseack; // @[MSHR.scala 186:28:chipyard.TestHarness.RocketConfig.fir@89355.4]
  assign io_schedule_bits_dir_valid = _T_77 | _T_91; // @[MSHR.scala 187:30:chipyard.TestHarness.RocketConfig.fir@89361.4]
  assign io_schedule_bits_dir_bits_set = request_set; // @[MSHR.scala 305:35:chipyard.TestHarness.RocketConfig.fir@89586.4]
  assign io_schedule_bits_dir_bits_way = meta_way; // @[MSHR.scala 306:35:chipyard.TestHarness.RocketConfig.fir@89587.4]
  assign io_schedule_bits_dir_bits_data_dirty = _T_76 ? 1'h0 : final_meta_writeback_dirty; // @[MSHR.scala 307:35:chipyard.TestHarness.RocketConfig.fir@89593.4]
  assign io_schedule_bits_dir_bits_data_state = _T_76 ? 2'h0 : final_meta_writeback_state; // @[MSHR.scala 307:35:chipyard.TestHarness.RocketConfig.fir@89593.4]
  assign io_schedule_bits_dir_bits_data_clients = _T_76 ? 1'h0 : final_meta_writeback_clients; // @[MSHR.scala 307:35:chipyard.TestHarness.RocketConfig.fir@89593.4]
  assign io_schedule_bits_dir_bits_data_tag = _T_76 ? 12'h0 : final_meta_writeback_tag; // @[MSHR.scala 307:35:chipyard.TestHarness.RocketConfig.fir@89593.4]
  assign io_schedule_bits_reload = _T_69 & w_grantack; // @[MSHR.scala 188:27:chipyard.TestHarness.RocketConfig.fir@89362.4]
  assign _GEN_170 = meta_valid & _T; // @[MSHR.scala 102:14:chipyard.TestHarness.RocketConfig.fir@89185.10]
  assign _GEN_174 = meta_valid & _T_10; // @[MSHR.scala 106:14:chipyard.TestHarness.RocketConfig.fir@89204.10]
  assign _GEN_176 = meta_valid & _T_15; // @[MSHR.scala 109:14:chipyard.TestHarness.RocketConfig.fir@89215.10]
  assign _GEN_180 = bad_grant & meta_hit; // @[MSHR.scala 251:14:chipyard.TestHarness.RocketConfig.fir@89498.10]
  assign _GEN_182 = _T_814 & new_request_prio_2; // @[MSHR.scala 582:14:chipyard.TestHarness.RocketConfig.fir@90634.10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  request_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  request_prio_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  request_prio_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  request_prio_2 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  request_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  request_opcode = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  request_param = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  request_size = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  request_source = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  request_tag = _RAND_9[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  request_offset = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  request_put = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  request_set = _RAND_12[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  meta_valid = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  meta_dirty = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  meta_state = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  meta_clients = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  meta_tag = _RAND_17[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  meta_hit = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  meta_way = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  s_rprobe = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  w_rprobeackfirst = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  w_rprobeacklast = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  s_release = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  w_releaseack = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  s_pprobe = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  s_acquire = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  s_flush = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  w_grantfirst = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  w_grantlast = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  w_grant = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  w_pprobeackfirst = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  w_pprobeacklast = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  w_pprobeack = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  s_grantack = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  s_execute = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  w_grantack = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  s_writeback = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  sink = _RAND_38[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  gotT = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  bad_grant = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  probes_done = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  probes_toN = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      request_valid <= 1'h0;
    end else begin
      request_valid <= _GEN_94;
    end
    if (io_allocate_valid) begin
      request_prio_0 <= io_allocate_bits_prio_0;
    end
    if (io_allocate_valid) begin
      request_prio_1 <= io_allocate_bits_prio_1;
    end
    if (io_allocate_valid) begin
      request_prio_2 <= io_allocate_bits_prio_2;
    end
    if (io_allocate_valid) begin
      request_control <= io_allocate_bits_control;
    end
    if (io_allocate_valid) begin
      request_opcode <= io_allocate_bits_opcode;
    end
    if (io_allocate_valid) begin
      request_param <= io_allocate_bits_param;
    end
    if (io_allocate_valid) begin
      request_size <= io_allocate_bits_size;
    end
    if (io_allocate_valid) begin
      request_source <= io_allocate_bits_source;
    end
    if (io_allocate_valid) begin
      request_tag <= io_allocate_bits_tag;
    end
    if (io_allocate_valid) begin
      request_offset <= io_allocate_bits_offset;
    end
    if (io_allocate_valid) begin
      request_put <= io_allocate_bits_put;
    end
    if (io_allocate_valid) begin
      request_set <= io_allocate_bits_set;
    end
    if (reset) begin
      meta_valid <= 1'h0;
    end else begin
      meta_valid <= _GEN_138;
    end
    if (_T_814) begin
      if (_T_760) begin
        if (bad_grant) begin
          meta_dirty <= 1'h0;
        end else if (request_prio_2) begin
          meta_dirty <= _T_120;
        end else if (request_control) begin
          if (meta_hit) begin
            meta_dirty <= 1'h0;
          end
        end else begin
          meta_dirty <= _T_139;
        end
      end else begin
        meta_dirty <= io_directory_bits_dirty;
      end
    end else if (io_sinkc_valid) begin
      meta_dirty <= _GEN_63;
    end else if (_T_33) begin
      meta_dirty <= _GEN_1;
    end
    if (_T_814) begin
      if (_T_760) begin
        if (bad_grant) begin
          if (meta_hit) begin
            meta_state <= 2'h1;
          end else begin
            meta_state <= 2'h0;
          end
        end else if (request_prio_2) begin
          if (_T_123) begin
            meta_state <= 2'h3;
          end
        end else if (request_control) begin
          if (meta_hit) begin
            meta_state <= 2'h0;
          end
        end else if (req_needT) begin
          if (_T_109) begin
            meta_state <= 2'h2;
          end else begin
            meta_state <= 2'h3;
          end
        end else if (_T_141) begin
          if (gotT) begin
            if (_T_109) begin
              meta_state <= 2'h2;
            end else begin
              meta_state <= 2'h3;
            end
          end else begin
            meta_state <= 2'h1;
          end
        end else if (_T_150) begin
          if (_T_144) begin
            meta_state <= 2'h2;
          end else begin
            meta_state <= 2'h3;
          end
        end else if (_T_148) begin
          meta_state <= 2'h3;
        end else begin
          meta_state <= 2'h1;
        end
      end else begin
        meta_state <= io_directory_bits_state;
      end
    end else if (_T_33) begin
      if (io_nestedwb_b_toB) begin
        meta_state <= 2'h1;
      end
    end
    if (_T_814) begin
      if (_T_760) begin
        if (bad_grant) begin
          meta_clients <= _T_156;
        end else if (request_prio_2) begin
          meta_clients <= _T_132;
        end else if (request_control) begin
          if (meta_hit) begin
            meta_clients <= _T_135;
          end
        end else begin
          meta_clients <= _T_158;
        end
      end else begin
        meta_clients <= io_directory_bits_clients;
      end
    end
    if (_T_814) begin
      if (_T_760) begin
        if (!(request_prio_2)) begin
          if (!(request_control)) begin
            meta_tag <= request_tag;
          end
        end
      end else begin
        meta_tag <= io_directory_bits_tag;
      end
    end
    if (_T_814) begin
      if (_T_760) begin
        if (!(bad_grant)) begin
          meta_hit <= _GEN_38;
        end
      end else begin
        meta_hit <= io_directory_bits_hit;
      end
    end else if (_T_33) begin
      if (io_nestedwb_b_toN) begin
        meta_hit <= 1'h0;
      end
    end
    if (_T_814) begin
      if (!(_T_760)) begin
        meta_way <= io_directory_bits_way;
      end
    end
    s_rprobe <= reset | _GEN_150;
    w_rprobeackfirst <= reset | _GEN_151;
    w_rprobeacklast <= reset | _GEN_152;
    s_release <= reset | _GEN_153;
    w_releaseack <= reset | _GEN_154;
    s_pprobe <= reset | _GEN_155;
    s_acquire <= reset | _GEN_156;
    s_flush <= reset | _GEN_157;
    w_grantfirst <= reset | _GEN_158;
    w_grantlast <= reset | _GEN_159;
    w_grant <= reset | _GEN_160;
    w_pprobeackfirst <= reset | _GEN_161;
    w_pprobeacklast <= reset | _GEN_162;
    w_pprobeack <= reset | _GEN_163;
    s_grantack <= reset | _GEN_165;
    s_execute <= reset | _GEN_166;
    w_grantack <= reset | _GEN_167;
    s_writeback <= reset | _GEN_168;
    if (io_sinkd_valid) begin
      if (_T_749) begin
        sink <= io_sinkd_bits_sink;
      end
    end
    if (_T_814) begin
      gotT <= 1'h0;
    end else if (io_sinkd_valid) begin
      if (_T_749) begin
        gotT <= _T_758;
      end
    end
    if (_T_814) begin
      bad_grant <= 1'h0;
    end else if (io_sinkd_valid) begin
      if (_T_749) begin
        bad_grant <= io_sinkd_bits_denied;
      end
    end
    if (_T_814) begin
      probes_done <= 1'h0;
    end else if (io_sinkc_valid) begin
      probes_done <= _T_713;
    end
    if (_T_814) begin
      probes_toN <= 1'h0;
    end else if (io_sinkc_valid) begin
      probes_toN <= _T_727;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_5) begin
          $fwrite(32'h80000002,"Assertion failed\n    at MSHR.scala:102 assert (!meta.clients.orR)\n"); // @[MSHR.scala 102:14:chipyard.TestHarness.RocketConfig.fir@89185.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_5) begin
          $fatal; // @[MSHR.scala 102:14:chipyard.TestHarness.RocketConfig.fir@89186.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_9) begin
          $fwrite(32'h80000002,"Assertion failed\n    at MSHR.scala:103 assert (!meta.dirty)\n"); // @[MSHR.scala 103:14:chipyard.TestHarness.RocketConfig.fir@89193.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_9) begin
          $fatal; // @[MSHR.scala 103:14:chipyard.TestHarness.RocketConfig.fir@89194.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_174 & _T_9) begin
          $fwrite(32'h80000002,"Assertion failed\n    at MSHR.scala:106 assert (!meta.dirty)\n"); // @[MSHR.scala 106:14:chipyard.TestHarness.RocketConfig.fir@89204.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_174 & _T_9) begin
          $fatal; // @[MSHR.scala 106:14:chipyard.TestHarness.RocketConfig.fir@89205.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_19) begin
          $fwrite(32'h80000002,"Assertion failed\n    at MSHR.scala:109 assert (meta.clients.orR)\n"); // @[MSHR.scala 109:14:chipyard.TestHarness.RocketConfig.fir@89215.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_19) begin
          $fatal; // @[MSHR.scala 109:14:chipyard.TestHarness.RocketConfig.fir@89216.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_26) begin
          $fwrite(32'h80000002,"Assertion failed\n    at MSHR.scala:110 assert ((meta.clients & (meta.clients - UInt(1))) === UInt(0)) // at most one\n"); // @[MSHR.scala 110:14:chipyard.TestHarness.RocketConfig.fir@89226.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_26) begin
          $fatal; // @[MSHR.scala 110:14:chipyard.TestHarness.RocketConfig.fir@89227.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_60) begin
          $fwrite(32'h80000002,"Assertion failed\n    at MSHR.scala:176 assert (!io.status.bits.nestB || !io.status.bits.blockB)\n"); // @[MSHR.scala 176:10:chipyard.TestHarness.RocketConfig.fir@89315.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_60) begin
          $fatal; // @[MSHR.scala 176:10:chipyard.TestHarness.RocketConfig.fir@89316.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_66) begin
          $fwrite(32'h80000002,"Assertion failed\n    at MSHR.scala:177 assert (!io.status.bits.nestC || !io.status.bits.blockC)\n"); // @[MSHR.scala 177:10:chipyard.TestHarness.RocketConfig.fir@89325.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_66) begin
          $fatal; // @[MSHR.scala 177:10:chipyard.TestHarness.RocketConfig.fir@89326.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_180 & _T_164) begin
          $fwrite(32'h80000002,"Assertion failed\n    at MSHR.scala:251 assert (!meta_valid || meta.state === BRANCH)\n"); // @[MSHR.scala 251:14:chipyard.TestHarness.RocketConfig.fir@89498.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_180 & _T_164) begin
          $fatal; // @[MSHR.scala 251:14:chipyard.TestHarness.RocketConfig.fir@89499.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_245 & _T_250) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH to evicted should be impossible (false,true,true,false,true)\n    at MSHR.scala:343 assert(!(evict === from.code), s\"State transition from ${from} to evicted should be impossible ${cfg}\")\n"); // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89698.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_245 & _T_250) begin
          $fatal; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89699.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_245 & _T_255) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH to flushed should be impossible (false,true,true,false,true)\n    at MSHR.scala:348 assert(!(before === from.code), s\"State transition from ${from} to flushed should be impossible ${cfg}\")\n"); // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89707.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_245 & _T_255) begin
          $fatal; // @[MSHR.scala 361:13:chipyard.TestHarness.RocketConfig.fir@89708.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_245 & _T_260) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH_C to evicted should be impossible (false,true,true,false,true)\n    at MSHR.scala:343 assert(!(evict === from.code), s\"State transition from ${from} to evicted should be impossible ${cfg}\")\n"); // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89716.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_245 & _T_260) begin
          $fatal; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89717.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_245 & _T_265) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH_C to flushed should be impossible (false,true,true,false,true)\n    at MSHR.scala:348 assert(!(before === from.code), s\"State transition from ${from} to flushed should be impossible ${cfg}\")\n"); // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89725.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_245 & _T_265) begin
          $fatal; // @[MSHR.scala 362:13:chipyard.TestHarness.RocketConfig.fir@89726.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_287) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_INVALID to S_BRANCH should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89753.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_287) begin
          $fatal; // @[MSHR.scala 372:15:chipyard.TestHarness.RocketConfig.fir@89754.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_294) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_INVALID to S_BRANCH_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 373:15:chipyard.TestHarness.RocketConfig.fir@89764.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_294) begin
          $fatal; // @[MSHR.scala 373:15:chipyard.TestHarness.RocketConfig.fir@89765.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_304) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_INVALID to S_TIP_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 375:15:chipyard.TestHarness.RocketConfig.fir@89778.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_304) begin
          $fatal; // @[MSHR.scala 375:15:chipyard.TestHarness.RocketConfig.fir@89779.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_311) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_INVALID to S_TIP_CD should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 376:15:chipyard.TestHarness.RocketConfig.fir@89789.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_311) begin
          $fatal; // @[MSHR.scala 376:15:chipyard.TestHarness.RocketConfig.fir@89790.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_324) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_INVALID to S_TRUNK_CD should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 379:15:chipyard.TestHarness.RocketConfig.fir@89806.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_324) begin
          $fatal; // @[MSHR.scala 379:15:chipyard.TestHarness.RocketConfig.fir@89807.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH to S_INVALID should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 381:15:chipyard.TestHarness.RocketConfig.fir@89817.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_331) begin
          $fatal; // @[MSHR.scala 381:15:chipyard.TestHarness.RocketConfig.fir@89818.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_338) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH to S_BRANCH_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 382:15:chipyard.TestHarness.RocketConfig.fir@89828.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_338) begin
          $fatal; // @[MSHR.scala 382:15:chipyard.TestHarness.RocketConfig.fir@89829.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_345) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH to S_TIP should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 383:15:chipyard.TestHarness.RocketConfig.fir@89839.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_345) begin
          $fatal; // @[MSHR.scala 383:15:chipyard.TestHarness.RocketConfig.fir@89840.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_352) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH to S_TIP_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 384:15:chipyard.TestHarness.RocketConfig.fir@89850.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_352) begin
          $fatal; // @[MSHR.scala 384:15:chipyard.TestHarness.RocketConfig.fir@89851.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_359) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH to S_TIP_CD should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 385:15:chipyard.TestHarness.RocketConfig.fir@89861.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_359) begin
          $fatal; // @[MSHR.scala 385:15:chipyard.TestHarness.RocketConfig.fir@89862.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_366) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH to S_TIP_D should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 386:15:chipyard.TestHarness.RocketConfig.fir@89872.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_366) begin
          $fatal; // @[MSHR.scala 386:15:chipyard.TestHarness.RocketConfig.fir@89873.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_373) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH to S_TRUNK_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 387:15:chipyard.TestHarness.RocketConfig.fir@89883.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_373) begin
          $fatal; // @[MSHR.scala 387:15:chipyard.TestHarness.RocketConfig.fir@89884.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_380) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH to S_TRUNK_CD should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 388:15:chipyard.TestHarness.RocketConfig.fir@89894.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_380) begin
          $fatal; // @[MSHR.scala 388:15:chipyard.TestHarness.RocketConfig.fir@89895.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_387) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH_C to S_INVALID should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 390:15:chipyard.TestHarness.RocketConfig.fir@89905.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_387) begin
          $fatal; // @[MSHR.scala 390:15:chipyard.TestHarness.RocketConfig.fir@89906.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_394) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH_C to S_BRANCH should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 391:15:chipyard.TestHarness.RocketConfig.fir@89916.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_394) begin
          $fatal; // @[MSHR.scala 391:15:chipyard.TestHarness.RocketConfig.fir@89917.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_401) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH_C to S_TIP should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 392:15:chipyard.TestHarness.RocketConfig.fir@89927.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_401) begin
          $fatal; // @[MSHR.scala 392:15:chipyard.TestHarness.RocketConfig.fir@89928.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_408) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH_C to S_TIP_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 393:15:chipyard.TestHarness.RocketConfig.fir@89938.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_408) begin
          $fatal; // @[MSHR.scala 393:15:chipyard.TestHarness.RocketConfig.fir@89939.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_415) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH_C to S_TIP_D should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 394:15:chipyard.TestHarness.RocketConfig.fir@89949.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_415) begin
          $fatal; // @[MSHR.scala 394:15:chipyard.TestHarness.RocketConfig.fir@89950.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_422) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH_C to S_TIP_CD should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 395:15:chipyard.TestHarness.RocketConfig.fir@89960.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_422) begin
          $fatal; // @[MSHR.scala 395:15:chipyard.TestHarness.RocketConfig.fir@89961.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_429) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH_C to S_TRUNK_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 396:15:chipyard.TestHarness.RocketConfig.fir@89971.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_429) begin
          $fatal; // @[MSHR.scala 396:15:chipyard.TestHarness.RocketConfig.fir@89972.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_436) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_BRANCH_C to S_TRUNK_CD should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 397:15:chipyard.TestHarness.RocketConfig.fir@89982.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_436) begin
          $fatal; // @[MSHR.scala 397:15:chipyard.TestHarness.RocketConfig.fir@89983.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_443) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP to S_INVALID should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 399:15:chipyard.TestHarness.RocketConfig.fir@89993.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_443) begin
          $fatal; // @[MSHR.scala 399:15:chipyard.TestHarness.RocketConfig.fir@89994.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_450) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP to S_BRANCH should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 400:15:chipyard.TestHarness.RocketConfig.fir@90004.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_450) begin
          $fatal; // @[MSHR.scala 400:15:chipyard.TestHarness.RocketConfig.fir@90005.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_457) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP to S_BRANCH_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 401:15:chipyard.TestHarness.RocketConfig.fir@90015.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_457) begin
          $fatal; // @[MSHR.scala 401:15:chipyard.TestHarness.RocketConfig.fir@90016.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_464) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP to S_TIP_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 402:15:chipyard.TestHarness.RocketConfig.fir@90026.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_464) begin
          $fatal; // @[MSHR.scala 402:15:chipyard.TestHarness.RocketConfig.fir@90027.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_474) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP to S_TIP_CD should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 404:15:chipyard.TestHarness.RocketConfig.fir@90040.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_474) begin
          $fatal; // @[MSHR.scala 404:15:chipyard.TestHarness.RocketConfig.fir@90041.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_484) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP to S_TRUNK_CD should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 406:15:chipyard.TestHarness.RocketConfig.fir@90054.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_484) begin
          $fatal; // @[MSHR.scala 406:15:chipyard.TestHarness.RocketConfig.fir@90055.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_491) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_C to S_INVALID should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 408:15:chipyard.TestHarness.RocketConfig.fir@90065.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_491) begin
          $fatal; // @[MSHR.scala 408:15:chipyard.TestHarness.RocketConfig.fir@90066.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_498) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_C to S_BRANCH should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 409:15:chipyard.TestHarness.RocketConfig.fir@90076.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_498) begin
          $fatal; // @[MSHR.scala 409:15:chipyard.TestHarness.RocketConfig.fir@90077.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_505) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_C to S_BRANCH_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 410:15:chipyard.TestHarness.RocketConfig.fir@90087.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_505) begin
          $fatal; // @[MSHR.scala 410:15:chipyard.TestHarness.RocketConfig.fir@90088.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_518) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_C to S_TIP_CD should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 413:15:chipyard.TestHarness.RocketConfig.fir@90104.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_518) begin
          $fatal; // @[MSHR.scala 413:15:chipyard.TestHarness.RocketConfig.fir@90105.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_528) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_C to S_TRUNK_CD should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 415:15:chipyard.TestHarness.RocketConfig.fir@90118.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_528) begin
          $fatal; // @[MSHR.scala 415:15:chipyard.TestHarness.RocketConfig.fir@90119.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_535) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_D to S_INVALID should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 417:15:chipyard.TestHarness.RocketConfig.fir@90129.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_535) begin
          $fatal; // @[MSHR.scala 417:15:chipyard.TestHarness.RocketConfig.fir@90130.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_542) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_D to S_BRANCH should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 418:15:chipyard.TestHarness.RocketConfig.fir@90140.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_542) begin
          $fatal; // @[MSHR.scala 418:15:chipyard.TestHarness.RocketConfig.fir@90141.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_549) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_D to S_BRANCH_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 419:15:chipyard.TestHarness.RocketConfig.fir@90151.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_549) begin
          $fatal; // @[MSHR.scala 419:15:chipyard.TestHarness.RocketConfig.fir@90152.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_556) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_D to S_TIP should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 420:15:chipyard.TestHarness.RocketConfig.fir@90162.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_556) begin
          $fatal; // @[MSHR.scala 420:15:chipyard.TestHarness.RocketConfig.fir@90163.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_563) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_D to S_TIP_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 421:15:chipyard.TestHarness.RocketConfig.fir@90173.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_563) begin
          $fatal; // @[MSHR.scala 421:15:chipyard.TestHarness.RocketConfig.fir@90174.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_570) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_D to S_TIP_CD should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 422:15:chipyard.TestHarness.RocketConfig.fir@90184.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_570) begin
          $fatal; // @[MSHR.scala 422:15:chipyard.TestHarness.RocketConfig.fir@90185.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_577) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_D to S_TRUNK_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 423:15:chipyard.TestHarness.RocketConfig.fir@90195.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_577) begin
          $fatal; // @[MSHR.scala 423:15:chipyard.TestHarness.RocketConfig.fir@90196.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_587) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_CD to S_INVALID should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 426:15:chipyard.TestHarness.RocketConfig.fir@90209.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_587) begin
          $fatal; // @[MSHR.scala 426:15:chipyard.TestHarness.RocketConfig.fir@90210.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_594) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_CD to S_BRANCH should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 427:15:chipyard.TestHarness.RocketConfig.fir@90220.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_594) begin
          $fatal; // @[MSHR.scala 427:15:chipyard.TestHarness.RocketConfig.fir@90221.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_601) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_CD to S_BRANCH_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 428:15:chipyard.TestHarness.RocketConfig.fir@90231.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_601) begin
          $fatal; // @[MSHR.scala 428:15:chipyard.TestHarness.RocketConfig.fir@90232.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_608) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_CD to S_TIP should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 429:15:chipyard.TestHarness.RocketConfig.fir@90242.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_608) begin
          $fatal; // @[MSHR.scala 429:15:chipyard.TestHarness.RocketConfig.fir@90243.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_615) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_CD to S_TIP_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 430:15:chipyard.TestHarness.RocketConfig.fir@90253.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_615) begin
          $fatal; // @[MSHR.scala 430:15:chipyard.TestHarness.RocketConfig.fir@90254.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_625) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TIP_CD to S_TRUNK_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 432:15:chipyard.TestHarness.RocketConfig.fir@90267.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_625) begin
          $fatal; // @[MSHR.scala 432:15:chipyard.TestHarness.RocketConfig.fir@90268.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_635) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TRUNK_C to S_INVALID should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 435:15:chipyard.TestHarness.RocketConfig.fir@90281.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_635) begin
          $fatal; // @[MSHR.scala 435:15:chipyard.TestHarness.RocketConfig.fir@90282.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_642) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TRUNK_C to S_BRANCH should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 436:15:chipyard.TestHarness.RocketConfig.fir@90292.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_642) begin
          $fatal; // @[MSHR.scala 436:15:chipyard.TestHarness.RocketConfig.fir@90293.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_649) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TRUNK_C to S_BRANCH_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 437:15:chipyard.TestHarness.RocketConfig.fir@90303.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_649) begin
          $fatal; // @[MSHR.scala 437:15:chipyard.TestHarness.RocketConfig.fir@90304.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_671) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TRUNK_CD to S_INVALID should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 444:15:chipyard.TestHarness.RocketConfig.fir@90329.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_671) begin
          $fatal; // @[MSHR.scala 444:15:chipyard.TestHarness.RocketConfig.fir@90330.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_678) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TRUNK_CD to S_BRANCH should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 445:15:chipyard.TestHarness.RocketConfig.fir@90340.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_678) begin
          $fatal; // @[MSHR.scala 445:15:chipyard.TestHarness.RocketConfig.fir@90341.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_685) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TRUNK_CD to S_BRANCH_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 446:15:chipyard.TestHarness.RocketConfig.fir@90351.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_685) begin
          $fatal; // @[MSHR.scala 446:15:chipyard.TestHarness.RocketConfig.fir@90352.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_692) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TRUNK_CD to S_TIP should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 447:15:chipyard.TestHarness.RocketConfig.fir@90362.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_692) begin
          $fatal; // @[MSHR.scala 447:15:chipyard.TestHarness.RocketConfig.fir@90363.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_699) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TRUNK_CD to S_TIP_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 448:15:chipyard.TestHarness.RocketConfig.fir@90373.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_699) begin
          $fatal; // @[MSHR.scala 448:15:chipyard.TestHarness.RocketConfig.fir@90374.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_280 & _T_712) begin
          $fwrite(32'h80000002,"Assertion failed: State transition from S_TRUNK_CD to S_TRUNK_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:356 assert(!(before === from.code && after === to.code), s\"State transition from ${from} to ${to} should be impossible ${cfg}\")\n"); // @[MSHR.scala 451:15:chipyard.TestHarness.RocketConfig.fir@90390.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_280 & _T_712) begin
          $fatal; // @[MSHR.scala 451:15:chipyard.TestHarness.RocketConfig.fir@90391.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_760 & _T_794) begin
          $fwrite(32'h80000002,"Assertion failed: State bypass from S_BRANCH should be impossible (false,true,true,false,true)\n    at MSHR.scala:513 assert(!(prior === from.code), s\"State bypass from ${from} should be impossible ${cfg}\")\n"); // @[MSHR.scala 519:11:chipyard.TestHarness.RocketConfig.fir@90539.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_760 & _T_794) begin
          $fatal; // @[MSHR.scala 519:11:chipyard.TestHarness.RocketConfig.fir@90540.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_760 & _T_799) begin
          $fwrite(32'h80000002,"Assertion failed: State bypass from S_BRANCH_C should be impossible (false,true,true,false,true)\n    at MSHR.scala:513 assert(!(prior === from.code), s\"State bypass from ${from} should be impossible ${cfg}\")\n"); // @[MSHR.scala 520:11:chipyard.TestHarness.RocketConfig.fir@90548.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_760 & _T_799) begin
          $fatal; // @[MSHR.scala 520:11:chipyard.TestHarness.RocketConfig.fir@90549.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_allocate_valid & _T_812) begin
          $fwrite(32'h80000002,"Assertion failed\n    at MSHR.scala:530 assert (!request_valid || (no_wait && io.schedule.fire()))\n"); // @[MSHR.scala 530:12:chipyard.TestHarness.RocketConfig.fir@90567.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_allocate_valid & _T_812) begin
          $fatal; // @[MSHR.scala 530:12:chipyard.TestHarness.RocketConfig.fir@90568.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_182 & _T_834) begin
          $fwrite(32'h80000002,"Assertion failed\n    at MSHR.scala:582 assert (new_meta.hit)\n"); // @[MSHR.scala 582:14:chipyard.TestHarness.RocketConfig.fir@90634.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_182 & _T_834) begin
          $fatal; // @[MSHR.scala 582:14:chipyard.TestHarness.RocketConfig.fir@90635.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
