module RoundAnyRawFNToRecFN_4( // @[:chipyard.TestHarness.RocketConfig.fir@237626.2]
  input         io_invalidExc, // @[:chipyard.TestHarness.RocketConfig.fir@237627.4]
  input         io_infiniteExc, // @[:chipyard.TestHarness.RocketConfig.fir@237627.4]
  input         io_in_isNaN, // @[:chipyard.TestHarness.RocketConfig.fir@237627.4]
  input         io_in_isInf, // @[:chipyard.TestHarness.RocketConfig.fir@237627.4]
  input         io_in_isZero, // @[:chipyard.TestHarness.RocketConfig.fir@237627.4]
  input         io_in_sign, // @[:chipyard.TestHarness.RocketConfig.fir@237627.4]
  input  [12:0] io_in_sExp, // @[:chipyard.TestHarness.RocketConfig.fir@237627.4]
  input  [55:0] io_in_sig, // @[:chipyard.TestHarness.RocketConfig.fir@237627.4]
  input  [2:0]  io_roundingMode, // @[:chipyard.TestHarness.RocketConfig.fir@237627.4]
  output [64:0] io_out, // @[:chipyard.TestHarness.RocketConfig.fir@237627.4]
  output [4:0]  io_exceptionFlags // @[:chipyard.TestHarness.RocketConfig.fir@237627.4]
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53:chipyard.TestHarness.RocketConfig.fir@237630.4]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53:chipyard.TestHarness.RocketConfig.fir@237632.4]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53:chipyard.TestHarness.RocketConfig.fir@237633.4]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53:chipyard.TestHarness.RocketConfig.fir@237634.4]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53:chipyard.TestHarness.RocketConfig.fir@237635.4]
  wire  _T; // @[RoundAnyRawFNToRecFN.scala 96:27:chipyard.TestHarness.RocketConfig.fir@237636.4]
  wire  _T_1; // @[RoundAnyRawFNToRecFN.scala 96:66:chipyard.TestHarness.RocketConfig.fir@237637.4]
  wire  _T_2; // @[RoundAnyRawFNToRecFN.scala 96:63:chipyard.TestHarness.RocketConfig.fir@237638.4]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42:chipyard.TestHarness.RocketConfig.fir@237639.4]
  wire  doShiftSigDown1; // @[RoundAnyRawFNToRecFN.scala 118:61:chipyard.TestHarness.RocketConfig.fir@237641.4]
  wire [11:0] _T_4; // @[primitives.scala 51:21:chipyard.TestHarness.RocketConfig.fir@237655.4]
  wire [64:0] _T_17; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@237668.4]
  wire [31:0] _T_23; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237674.4]
  wire [31:0] _T_25; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237676.4]
  wire [31:0] _T_27; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237678.4]
  wire [31:0] _T_28; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237679.4]
  wire [31:0] _GEN_0; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237684.4]
  wire [31:0] _T_33; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237684.4]
  wire [31:0] _T_35; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237686.4]
  wire [31:0] _T_37; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237688.4]
  wire [31:0] _T_38; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237689.4]
  wire [31:0] _GEN_1; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237694.4]
  wire [31:0] _T_43; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237694.4]
  wire [31:0] _T_45; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237696.4]
  wire [31:0] _T_47; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237698.4]
  wire [31:0] _T_48; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237699.4]
  wire [31:0] _GEN_2; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237704.4]
  wire [31:0] _T_53; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237704.4]
  wire [31:0] _T_55; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237706.4]
  wire [31:0] _T_57; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237708.4]
  wire [31:0] _T_58; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237709.4]
  wire [31:0] _GEN_3; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237714.4]
  wire [31:0] _T_63; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237714.4]
  wire [31:0] _T_65; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237716.4]
  wire [31:0] _T_67; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237718.4]
  wire [31:0] _T_68; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237719.4]
  wire [15:0] _T_74; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237725.4]
  wire [15:0] _T_76; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237727.4]
  wire [15:0] _T_78; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237729.4]
  wire [15:0] _T_79; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237730.4]
  wire [15:0] _GEN_4; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237735.4]
  wire [15:0] _T_84; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237735.4]
  wire [15:0] _T_86; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237737.4]
  wire [15:0] _T_88; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237739.4]
  wire [15:0] _T_89; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237740.4]
  wire [15:0] _GEN_5; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237745.4]
  wire [15:0] _T_94; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237745.4]
  wire [15:0] _T_96; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237747.4]
  wire [15:0] _T_98; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237749.4]
  wire [15:0] _T_99; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237750.4]
  wire [15:0] _GEN_6; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237755.4]
  wire [15:0] _T_104; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237755.4]
  wire [15:0] _T_106; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237757.4]
  wire [15:0] _T_108; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237759.4]
  wire [15:0] _T_109; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237760.4]
  wire [50:0] _T_118; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237769.4]
  wire [50:0] _T_119; // @[primitives.scala 74:36:chipyard.TestHarness.RocketConfig.fir@237770.4]
  wire [50:0] _T_120; // @[primitives.scala 74:21:chipyard.TestHarness.RocketConfig.fir@237771.4]
  wire [50:0] _T_121; // @[primitives.scala 74:17:chipyard.TestHarness.RocketConfig.fir@237772.4]
  wire [50:0] _T_122; // @[primitives.scala 74:36:chipyard.TestHarness.RocketConfig.fir@237773.4]
  wire [50:0] _T_123; // @[primitives.scala 74:21:chipyard.TestHarness.RocketConfig.fir@237774.4]
  wire [50:0] _T_124; // @[primitives.scala 74:17:chipyard.TestHarness.RocketConfig.fir@237775.4]
  wire [50:0] _T_125; // @[primitives.scala 74:36:chipyard.TestHarness.RocketConfig.fir@237776.4]
  wire [50:0] _T_126; // @[primitives.scala 74:21:chipyard.TestHarness.RocketConfig.fir@237777.4]
  wire [50:0] _T_127; // @[primitives.scala 74:17:chipyard.TestHarness.RocketConfig.fir@237778.4]
  wire [50:0] _T_128; // @[primitives.scala 74:36:chipyard.TestHarness.RocketConfig.fir@237779.4]
  wire [50:0] _T_129; // @[primitives.scala 74:21:chipyard.TestHarness.RocketConfig.fir@237780.4]
  wire [50:0] _T_130; // @[primitives.scala 74:17:chipyard.TestHarness.RocketConfig.fir@237781.4]
  wire [53:0] _T_131; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237782.4]
  wire [2:0] _T_147; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237798.4]
  wire [2:0] _T_148; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@237799.4]
  wire [2:0] _T_149; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@237800.4]
  wire [2:0] _T_150; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@237801.4]
  wire [2:0] _T_151; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@237802.4]
  wire [53:0] _T_152; // @[primitives.scala 66:24:chipyard.TestHarness.RocketConfig.fir@237803.4]
  wire [53:0] _T_153; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@237804.4]
  wire [53:0] _GEN_7; // @[RoundAnyRawFNToRecFN.scala 157:23:chipyard.TestHarness.RocketConfig.fir@237805.4]
  wire [53:0] _T_154; // @[RoundAnyRawFNToRecFN.scala 157:23:chipyard.TestHarness.RocketConfig.fir@237805.4]
  wire [55:0] _T_155; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237806.4]
  wire [55:0] _T_157; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237808.4]
  wire [55:0] _T_158; // @[RoundAnyRawFNToRecFN.scala 161:28:chipyard.TestHarness.RocketConfig.fir@237809.4]
  wire [55:0] _T_159; // @[RoundAnyRawFNToRecFN.scala 161:46:chipyard.TestHarness.RocketConfig.fir@237810.4]
  wire [55:0] _T_160; // @[RoundAnyRawFNToRecFN.scala 162:40:chipyard.TestHarness.RocketConfig.fir@237811.4]
  wire  _T_161; // @[RoundAnyRawFNToRecFN.scala 162:56:chipyard.TestHarness.RocketConfig.fir@237812.4]
  wire [55:0] _T_162; // @[RoundAnyRawFNToRecFN.scala 163:42:chipyard.TestHarness.RocketConfig.fir@237813.4]
  wire  _T_163; // @[RoundAnyRawFNToRecFN.scala 163:62:chipyard.TestHarness.RocketConfig.fir@237814.4]
  wire  _T_164; // @[RoundAnyRawFNToRecFN.scala 164:36:chipyard.TestHarness.RocketConfig.fir@237815.4]
  wire  _T_165; // @[RoundAnyRawFNToRecFN.scala 167:38:chipyard.TestHarness.RocketConfig.fir@237816.4]
  wire  _T_166; // @[RoundAnyRawFNToRecFN.scala 167:67:chipyard.TestHarness.RocketConfig.fir@237817.4]
  wire  _T_167; // @[RoundAnyRawFNToRecFN.scala 169:29:chipyard.TestHarness.RocketConfig.fir@237818.4]
  wire  _T_168; // @[RoundAnyRawFNToRecFN.scala 168:31:chipyard.TestHarness.RocketConfig.fir@237819.4]
  wire [55:0] _T_169; // @[RoundAnyRawFNToRecFN.scala 172:32:chipyard.TestHarness.RocketConfig.fir@237820.4]
  wire [54:0] _T_171; // @[RoundAnyRawFNToRecFN.scala 172:49:chipyard.TestHarness.RocketConfig.fir@237822.4]
  wire  _T_172; // @[RoundAnyRawFNToRecFN.scala 173:49:chipyard.TestHarness.RocketConfig.fir@237823.4]
  wire  _T_173; // @[RoundAnyRawFNToRecFN.scala 174:30:chipyard.TestHarness.RocketConfig.fir@237824.4]
  wire  _T_174; // @[RoundAnyRawFNToRecFN.scala 173:64:chipyard.TestHarness.RocketConfig.fir@237825.4]
  wire [54:0] _T_176; // @[RoundAnyRawFNToRecFN.scala 173:25:chipyard.TestHarness.RocketConfig.fir@237827.4]
  wire [54:0] _T_177; // @[RoundAnyRawFNToRecFN.scala 173:21:chipyard.TestHarness.RocketConfig.fir@237828.4]
  wire [54:0] _T_178; // @[RoundAnyRawFNToRecFN.scala 172:61:chipyard.TestHarness.RocketConfig.fir@237829.4]
  wire [55:0] _T_179; // @[RoundAnyRawFNToRecFN.scala 178:32:chipyard.TestHarness.RocketConfig.fir@237830.4]
  wire [55:0] _T_180; // @[RoundAnyRawFNToRecFN.scala 178:30:chipyard.TestHarness.RocketConfig.fir@237831.4]
  wire  _T_182; // @[RoundAnyRawFNToRecFN.scala 179:42:chipyard.TestHarness.RocketConfig.fir@237833.4]
  wire [54:0] _T_184; // @[RoundAnyRawFNToRecFN.scala 179:24:chipyard.TestHarness.RocketConfig.fir@237835.4]
  wire [54:0] _GEN_8; // @[RoundAnyRawFNToRecFN.scala 178:47:chipyard.TestHarness.RocketConfig.fir@237836.4]
  wire [54:0] _T_185; // @[RoundAnyRawFNToRecFN.scala 178:47:chipyard.TestHarness.RocketConfig.fir@237836.4]
  wire [54:0] _T_186; // @[RoundAnyRawFNToRecFN.scala 171:16:chipyard.TestHarness.RocketConfig.fir@237837.4]
  wire [2:0] _T_188; // @[RoundAnyRawFNToRecFN.scala 183:69:chipyard.TestHarness.RocketConfig.fir@237839.4]
  wire [12:0] _GEN_9; // @[RoundAnyRawFNToRecFN.scala 183:40:chipyard.TestHarness.RocketConfig.fir@237840.4]
  wire [13:0] _T_189; // @[RoundAnyRawFNToRecFN.scala 183:40:chipyard.TestHarness.RocketConfig.fir@237840.4]
  wire [11:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37:chipyard.TestHarness.RocketConfig.fir@237841.4]
  wire [51:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 187:16:chipyard.TestHarness.RocketConfig.fir@237845.4]
  wire [3:0] _T_194; // @[RoundAnyRawFNToRecFN.scala 194:30:chipyard.TestHarness.RocketConfig.fir@237847.4]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50:chipyard.TestHarness.RocketConfig.fir@237848.4]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31:chipyard.TestHarness.RocketConfig.fir@237850.4]
  wire  _T_199; // @[RoundAnyRawFNToRecFN.scala 201:16:chipyard.TestHarness.RocketConfig.fir@237854.4]
  wire  _T_201; // @[RoundAnyRawFNToRecFN.scala 203:30:chipyard.TestHarness.RocketConfig.fir@237856.4]
  wire  _T_203; // @[RoundAnyRawFNToRecFN.scala 203:70:chipyard.TestHarness.RocketConfig.fir@237858.4]
  wire  _T_204; // @[RoundAnyRawFNToRecFN.scala 203:49:chipyard.TestHarness.RocketConfig.fir@237859.4]
  wire  _T_206; // @[RoundAnyRawFNToRecFN.scala 205:67:chipyard.TestHarness.RocketConfig.fir@237861.4]
  wire  _T_207; // @[RoundAnyRawFNToRecFN.scala 207:29:chipyard.TestHarness.RocketConfig.fir@237862.4]
  wire  _T_208; // @[RoundAnyRawFNToRecFN.scala 206:46:chipyard.TestHarness.RocketConfig.fir@237863.4]
  wire  _T_211; // @[RoundAnyRawFNToRecFN.scala 209:16:chipyard.TestHarness.RocketConfig.fir@237866.4]
  wire [1:0] _T_212; // @[RoundAnyRawFNToRecFN.scala 218:48:chipyard.TestHarness.RocketConfig.fir@237867.4]
  wire  _T_213; // @[RoundAnyRawFNToRecFN.scala 218:62:chipyard.TestHarness.RocketConfig.fir@237868.4]
  wire  _T_214; // @[RoundAnyRawFNToRecFN.scala 218:32:chipyard.TestHarness.RocketConfig.fir@237869.4]
  wire  _T_217; // @[RoundAnyRawFNToRecFN.scala 219:30:chipyard.TestHarness.RocketConfig.fir@237872.4]
  wire  _T_218; // @[RoundAnyRawFNToRecFN.scala 218:74:chipyard.TestHarness.RocketConfig.fir@237873.4]
  wire  _T_222; // @[RoundAnyRawFNToRecFN.scala 221:39:chipyard.TestHarness.RocketConfig.fir@237877.4]
  wire  _T_223; // @[RoundAnyRawFNToRecFN.scala 221:34:chipyard.TestHarness.RocketConfig.fir@237878.4]
  wire  _T_225; // @[RoundAnyRawFNToRecFN.scala 224:38:chipyard.TestHarness.RocketConfig.fir@237880.4]
  wire  _T_226; // @[RoundAnyRawFNToRecFN.scala 225:45:chipyard.TestHarness.RocketConfig.fir@237881.4]
  wire  _T_227; // @[RoundAnyRawFNToRecFN.scala 225:60:chipyard.TestHarness.RocketConfig.fir@237882.4]
  wire  _T_228; // @[RoundAnyRawFNToRecFN.scala 220:27:chipyard.TestHarness.RocketConfig.fir@237883.4]
  wire  _T_229; // @[RoundAnyRawFNToRecFN.scala 219:76:chipyard.TestHarness.RocketConfig.fir@237884.4]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40:chipyard.TestHarness.RocketConfig.fir@237885.4]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49:chipyard.TestHarness.RocketConfig.fir@237887.4]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34:chipyard.TestHarness.RocketConfig.fir@237889.4]
  wire  notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 234:49:chipyard.TestHarness.RocketConfig.fir@237890.4]
  wire  _T_232; // @[RoundAnyRawFNToRecFN.scala 235:22:chipyard.TestHarness.RocketConfig.fir@237891.4]
  wire  _T_233; // @[RoundAnyRawFNToRecFN.scala 235:36:chipyard.TestHarness.RocketConfig.fir@237892.4]
  wire  _T_234; // @[RoundAnyRawFNToRecFN.scala 235:33:chipyard.TestHarness.RocketConfig.fir@237893.4]
  wire  _T_235; // @[RoundAnyRawFNToRecFN.scala 235:64:chipyard.TestHarness.RocketConfig.fir@237894.4]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61:chipyard.TestHarness.RocketConfig.fir@237895.4]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32:chipyard.TestHarness.RocketConfig.fir@237896.4]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32:chipyard.TestHarness.RocketConfig.fir@237897.4]
  wire  _T_236; // @[RoundAnyRawFNToRecFN.scala 238:43:chipyard.TestHarness.RocketConfig.fir@237898.4]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28:chipyard.TestHarness.RocketConfig.fir@237899.4]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60:chipyard.TestHarness.RocketConfig.fir@237901.4]
  wire  _T_238; // @[RoundAnyRawFNToRecFN.scala 243:20:chipyard.TestHarness.RocketConfig.fir@237902.4]
  wire  _T_239; // @[RoundAnyRawFNToRecFN.scala 243:60:chipyard.TestHarness.RocketConfig.fir@237903.4]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45:chipyard.TestHarness.RocketConfig.fir@237904.4]
  wire  _T_240; // @[RoundAnyRawFNToRecFN.scala 244:42:chipyard.TestHarness.RocketConfig.fir@237905.4]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39:chipyard.TestHarness.RocketConfig.fir@237906.4]
  wire  _T_241; // @[RoundAnyRawFNToRecFN.scala 246:45:chipyard.TestHarness.RocketConfig.fir@237907.4]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32:chipyard.TestHarness.RocketConfig.fir@237908.4]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22:chipyard.TestHarness.RocketConfig.fir@237909.4]
  wire  _T_242; // @[RoundAnyRawFNToRecFN.scala 251:32:chipyard.TestHarness.RocketConfig.fir@237910.4]
  wire [11:0] _T_243; // @[RoundAnyRawFNToRecFN.scala 251:18:chipyard.TestHarness.RocketConfig.fir@237911.4]
  wire [11:0] _T_244; // @[RoundAnyRawFNToRecFN.scala 251:14:chipyard.TestHarness.RocketConfig.fir@237912.4]
  wire [11:0] _T_245; // @[RoundAnyRawFNToRecFN.scala 250:24:chipyard.TestHarness.RocketConfig.fir@237913.4]
  wire [11:0] _T_247; // @[RoundAnyRawFNToRecFN.scala 255:18:chipyard.TestHarness.RocketConfig.fir@237915.4]
  wire [11:0] _T_248; // @[RoundAnyRawFNToRecFN.scala 255:14:chipyard.TestHarness.RocketConfig.fir@237916.4]
  wire [11:0] _T_249; // @[RoundAnyRawFNToRecFN.scala 254:17:chipyard.TestHarness.RocketConfig.fir@237917.4]
  wire [11:0] _T_250; // @[RoundAnyRawFNToRecFN.scala 259:18:chipyard.TestHarness.RocketConfig.fir@237918.4]
  wire [11:0] _T_251; // @[RoundAnyRawFNToRecFN.scala 259:14:chipyard.TestHarness.RocketConfig.fir@237919.4]
  wire [11:0] _T_252; // @[RoundAnyRawFNToRecFN.scala 258:17:chipyard.TestHarness.RocketConfig.fir@237920.4]
  wire [11:0] _T_253; // @[RoundAnyRawFNToRecFN.scala 263:18:chipyard.TestHarness.RocketConfig.fir@237921.4]
  wire [11:0] _T_254; // @[RoundAnyRawFNToRecFN.scala 263:14:chipyard.TestHarness.RocketConfig.fir@237922.4]
  wire [11:0] _T_255; // @[RoundAnyRawFNToRecFN.scala 262:17:chipyard.TestHarness.RocketConfig.fir@237923.4]
  wire [11:0] _T_256; // @[RoundAnyRawFNToRecFN.scala 267:16:chipyard.TestHarness.RocketConfig.fir@237924.4]
  wire [11:0] _T_257; // @[RoundAnyRawFNToRecFN.scala 266:18:chipyard.TestHarness.RocketConfig.fir@237925.4]
  wire [11:0] _T_258; // @[RoundAnyRawFNToRecFN.scala 271:16:chipyard.TestHarness.RocketConfig.fir@237926.4]
  wire [11:0] _T_259; // @[RoundAnyRawFNToRecFN.scala 270:15:chipyard.TestHarness.RocketConfig.fir@237927.4]
  wire [11:0] _T_260; // @[RoundAnyRawFNToRecFN.scala 275:16:chipyard.TestHarness.RocketConfig.fir@237928.4]
  wire [11:0] _T_261; // @[RoundAnyRawFNToRecFN.scala 274:15:chipyard.TestHarness.RocketConfig.fir@237929.4]
  wire [11:0] _T_262; // @[RoundAnyRawFNToRecFN.scala 276:16:chipyard.TestHarness.RocketConfig.fir@237930.4]
  wire [11:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77:chipyard.TestHarness.RocketConfig.fir@237931.4]
  wire  _T_263; // @[RoundAnyRawFNToRecFN.scala 278:22:chipyard.TestHarness.RocketConfig.fir@237932.4]
  wire  _T_264; // @[RoundAnyRawFNToRecFN.scala 278:38:chipyard.TestHarness.RocketConfig.fir@237933.4]
  wire [51:0] _T_265; // @[RoundAnyRawFNToRecFN.scala 279:16:chipyard.TestHarness.RocketConfig.fir@237934.4]
  wire [51:0] _T_266; // @[RoundAnyRawFNToRecFN.scala 278:12:chipyard.TestHarness.RocketConfig.fir@237935.4]
  wire [51:0] _T_268; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@237937.4]
  wire [51:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11:chipyard.TestHarness.RocketConfig.fir@237938.4]
  wire [12:0] _T_269; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237939.4]
  wire [1:0] _T_271; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237942.4]
  wire [2:0] _T_273; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237944.4]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53:chipyard.TestHarness.RocketConfig.fir@237630.4]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53:chipyard.TestHarness.RocketConfig.fir@237632.4]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53:chipyard.TestHarness.RocketConfig.fir@237633.4]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53:chipyard.TestHarness.RocketConfig.fir@237634.4]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53:chipyard.TestHarness.RocketConfig.fir@237635.4]
  assign _T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27:chipyard.TestHarness.RocketConfig.fir@237636.4]
  assign _T_1 = ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:66:chipyard.TestHarness.RocketConfig.fir@237637.4]
  assign _T_2 = roundingMode_max & _T_1; // @[RoundAnyRawFNToRecFN.scala 96:63:chipyard.TestHarness.RocketConfig.fir@237638.4]
  assign roundMagUp = _T | _T_2; // @[RoundAnyRawFNToRecFN.scala 96:42:chipyard.TestHarness.RocketConfig.fir@237639.4]
  assign doShiftSigDown1 = io_in_sig[55]; // @[RoundAnyRawFNToRecFN.scala 118:61:chipyard.TestHarness.RocketConfig.fir@237641.4]
  assign _T_4 = ~io_in_sExp[11:0]; // @[primitives.scala 51:21:chipyard.TestHarness.RocketConfig.fir@237655.4]
  assign _T_17 = -65'sh10000000000000000 >>> _T_4[5:0]; // @[primitives.scala 77:58:chipyard.TestHarness.RocketConfig.fir@237668.4]
  assign _T_23 = {{16'd0}, _T_17[44:29]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237674.4]
  assign _T_25 = {_T_17[28:13], 16'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237676.4]
  assign _T_27 = _T_25 & 32'hffff0000; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237678.4]
  assign _T_28 = _T_23 | _T_27; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237679.4]
  assign _GEN_0 = {{8'd0}, _T_28[31:8]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237684.4]
  assign _T_33 = _GEN_0 & 32'hff00ff; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237684.4]
  assign _T_35 = {_T_28[23:0], 8'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237686.4]
  assign _T_37 = _T_35 & 32'hff00ff00; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237688.4]
  assign _T_38 = _T_33 | _T_37; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237689.4]
  assign _GEN_1 = {{4'd0}, _T_38[31:4]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237694.4]
  assign _T_43 = _GEN_1 & 32'hf0f0f0f; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237694.4]
  assign _T_45 = {_T_38[27:0], 4'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237696.4]
  assign _T_47 = _T_45 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237698.4]
  assign _T_48 = _T_43 | _T_47; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237699.4]
  assign _GEN_2 = {{2'd0}, _T_48[31:2]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237704.4]
  assign _T_53 = _GEN_2 & 32'h33333333; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237704.4]
  assign _T_55 = {_T_48[29:0], 2'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237706.4]
  assign _T_57 = _T_55 & 32'hcccccccc; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237708.4]
  assign _T_58 = _T_53 | _T_57; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237709.4]
  assign _GEN_3 = {{1'd0}, _T_58[31:1]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237714.4]
  assign _T_63 = _GEN_3 & 32'h55555555; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237714.4]
  assign _T_65 = {_T_58[30:0], 1'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237716.4]
  assign _T_67 = _T_65 & 32'haaaaaaaa; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237718.4]
  assign _T_68 = _T_63 | _T_67; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237719.4]
  assign _T_74 = {{8'd0}, _T_17[60:53]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237725.4]
  assign _T_76 = {_T_17[52:45], 8'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237727.4]
  assign _T_78 = _T_76 & 16'hff00; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237729.4]
  assign _T_79 = _T_74 | _T_78; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237730.4]
  assign _GEN_4 = {{4'd0}, _T_79[15:4]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237735.4]
  assign _T_84 = _GEN_4 & 16'hf0f; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237735.4]
  assign _T_86 = {_T_79[11:0], 4'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237737.4]
  assign _T_88 = _T_86 & 16'hf0f0; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237739.4]
  assign _T_89 = _T_84 | _T_88; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237740.4]
  assign _GEN_5 = {{2'd0}, _T_89[15:2]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237745.4]
  assign _T_94 = _GEN_5 & 16'h3333; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237745.4]
  assign _T_96 = {_T_89[13:0], 2'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237747.4]
  assign _T_98 = _T_96 & 16'hcccc; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237749.4]
  assign _T_99 = _T_94 | _T_98; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237750.4]
  assign _GEN_6 = {{1'd0}, _T_99[15:1]}; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237755.4]
  assign _T_104 = _GEN_6 & 16'h5555; // @[Bitwise.scala 103:31:chipyard.TestHarness.RocketConfig.fir@237755.4]
  assign _T_106 = {_T_99[14:0], 1'h0}; // @[Bitwise.scala 103:65:chipyard.TestHarness.RocketConfig.fir@237757.4]
  assign _T_108 = _T_106 & 16'haaaa; // @[Bitwise.scala 103:75:chipyard.TestHarness.RocketConfig.fir@237759.4]
  assign _T_109 = _T_104 | _T_108; // @[Bitwise.scala 103:39:chipyard.TestHarness.RocketConfig.fir@237760.4]
  assign _T_118 = {_T_68,_T_109,_T_17[61],_T_17[62],_T_17[63]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237769.4]
  assign _T_119 = ~_T_118; // @[primitives.scala 74:36:chipyard.TestHarness.RocketConfig.fir@237770.4]
  assign _T_120 = _T_4[6] ? 51'h0 : _T_119; // @[primitives.scala 74:21:chipyard.TestHarness.RocketConfig.fir@237771.4]
  assign _T_121 = ~_T_120; // @[primitives.scala 74:17:chipyard.TestHarness.RocketConfig.fir@237772.4]
  assign _T_122 = ~_T_121; // @[primitives.scala 74:36:chipyard.TestHarness.RocketConfig.fir@237773.4]
  assign _T_123 = _T_4[7] ? 51'h0 : _T_122; // @[primitives.scala 74:21:chipyard.TestHarness.RocketConfig.fir@237774.4]
  assign _T_124 = ~_T_123; // @[primitives.scala 74:17:chipyard.TestHarness.RocketConfig.fir@237775.4]
  assign _T_125 = ~_T_124; // @[primitives.scala 74:36:chipyard.TestHarness.RocketConfig.fir@237776.4]
  assign _T_126 = _T_4[8] ? 51'h0 : _T_125; // @[primitives.scala 74:21:chipyard.TestHarness.RocketConfig.fir@237777.4]
  assign _T_127 = ~_T_126; // @[primitives.scala 74:17:chipyard.TestHarness.RocketConfig.fir@237778.4]
  assign _T_128 = ~_T_127; // @[primitives.scala 74:36:chipyard.TestHarness.RocketConfig.fir@237779.4]
  assign _T_129 = _T_4[9] ? 51'h0 : _T_128; // @[primitives.scala 74:21:chipyard.TestHarness.RocketConfig.fir@237780.4]
  assign _T_130 = ~_T_129; // @[primitives.scala 74:17:chipyard.TestHarness.RocketConfig.fir@237781.4]
  assign _T_131 = {_T_130,3'h7}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237782.4]
  assign _T_147 = {_T_17[0],_T_17[1],_T_17[2]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237798.4]
  assign _T_148 = _T_4[6] ? _T_147 : 3'h0; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@237799.4]
  assign _T_149 = _T_4[7] ? _T_148 : 3'h0; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@237800.4]
  assign _T_150 = _T_4[8] ? _T_149 : 3'h0; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@237801.4]
  assign _T_151 = _T_4[9] ? _T_150 : 3'h0; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@237802.4]
  assign _T_152 = _T_4[10] ? _T_131 : {{51'd0}, _T_151}; // @[primitives.scala 66:24:chipyard.TestHarness.RocketConfig.fir@237803.4]
  assign _T_153 = _T_4[11] ? _T_152 : 54'h0; // @[primitives.scala 61:24:chipyard.TestHarness.RocketConfig.fir@237804.4]
  assign _GEN_7 = {{53'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23:chipyard.TestHarness.RocketConfig.fir@237805.4]
  assign _T_154 = _T_153 | _GEN_7; // @[RoundAnyRawFNToRecFN.scala 157:23:chipyard.TestHarness.RocketConfig.fir@237805.4]
  assign _T_155 = {_T_154,2'h3}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237806.4]
  assign _T_157 = {1'h0,_T_155[55:1]}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237808.4]
  assign _T_158 = ~_T_157; // @[RoundAnyRawFNToRecFN.scala 161:28:chipyard.TestHarness.RocketConfig.fir@237809.4]
  assign _T_159 = _T_158 & _T_155; // @[RoundAnyRawFNToRecFN.scala 161:46:chipyard.TestHarness.RocketConfig.fir@237810.4]
  assign _T_160 = io_in_sig & _T_159; // @[RoundAnyRawFNToRecFN.scala 162:40:chipyard.TestHarness.RocketConfig.fir@237811.4]
  assign _T_161 = |_T_160; // @[RoundAnyRawFNToRecFN.scala 162:56:chipyard.TestHarness.RocketConfig.fir@237812.4]
  assign _T_162 = io_in_sig & _T_157; // @[RoundAnyRawFNToRecFN.scala 163:42:chipyard.TestHarness.RocketConfig.fir@237813.4]
  assign _T_163 = |_T_162; // @[RoundAnyRawFNToRecFN.scala 163:62:chipyard.TestHarness.RocketConfig.fir@237814.4]
  assign _T_164 = _T_161 | _T_163; // @[RoundAnyRawFNToRecFN.scala 164:36:chipyard.TestHarness.RocketConfig.fir@237815.4]
  assign _T_165 = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38:chipyard.TestHarness.RocketConfig.fir@237816.4]
  assign _T_166 = _T_165 & _T_161; // @[RoundAnyRawFNToRecFN.scala 167:67:chipyard.TestHarness.RocketConfig.fir@237817.4]
  assign _T_167 = roundMagUp & _T_164; // @[RoundAnyRawFNToRecFN.scala 169:29:chipyard.TestHarness.RocketConfig.fir@237818.4]
  assign _T_168 = _T_166 | _T_167; // @[RoundAnyRawFNToRecFN.scala 168:31:chipyard.TestHarness.RocketConfig.fir@237819.4]
  assign _T_169 = io_in_sig | _T_155; // @[RoundAnyRawFNToRecFN.scala 172:32:chipyard.TestHarness.RocketConfig.fir@237820.4]
  assign _T_171 = _T_169[55:2] + 54'h1; // @[RoundAnyRawFNToRecFN.scala 172:49:chipyard.TestHarness.RocketConfig.fir@237822.4]
  assign _T_172 = roundingMode_near_even & _T_161; // @[RoundAnyRawFNToRecFN.scala 173:49:chipyard.TestHarness.RocketConfig.fir@237823.4]
  assign _T_173 = ~_T_163; // @[RoundAnyRawFNToRecFN.scala 174:30:chipyard.TestHarness.RocketConfig.fir@237824.4]
  assign _T_174 = _T_172 & _T_173; // @[RoundAnyRawFNToRecFN.scala 173:64:chipyard.TestHarness.RocketConfig.fir@237825.4]
  assign _T_176 = _T_174 ? _T_155[55:1] : 55'h0; // @[RoundAnyRawFNToRecFN.scala 173:25:chipyard.TestHarness.RocketConfig.fir@237827.4]
  assign _T_177 = ~_T_176; // @[RoundAnyRawFNToRecFN.scala 173:21:chipyard.TestHarness.RocketConfig.fir@237828.4]
  assign _T_178 = _T_171 & _T_177; // @[RoundAnyRawFNToRecFN.scala 172:61:chipyard.TestHarness.RocketConfig.fir@237829.4]
  assign _T_179 = ~_T_155; // @[RoundAnyRawFNToRecFN.scala 178:32:chipyard.TestHarness.RocketConfig.fir@237830.4]
  assign _T_180 = io_in_sig & _T_179; // @[RoundAnyRawFNToRecFN.scala 178:30:chipyard.TestHarness.RocketConfig.fir@237831.4]
  assign _T_182 = roundingMode_odd & _T_164; // @[RoundAnyRawFNToRecFN.scala 179:42:chipyard.TestHarness.RocketConfig.fir@237833.4]
  assign _T_184 = _T_182 ? _T_159[55:1] : 55'h0; // @[RoundAnyRawFNToRecFN.scala 179:24:chipyard.TestHarness.RocketConfig.fir@237835.4]
  assign _GEN_8 = {{1'd0}, _T_180[55:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47:chipyard.TestHarness.RocketConfig.fir@237836.4]
  assign _T_185 = _GEN_8 | _T_184; // @[RoundAnyRawFNToRecFN.scala 178:47:chipyard.TestHarness.RocketConfig.fir@237836.4]
  assign _T_186 = _T_168 ? _T_178 : _T_185; // @[RoundAnyRawFNToRecFN.scala 171:16:chipyard.TestHarness.RocketConfig.fir@237837.4]
  assign _T_188 = {1'b0,$signed(_T_186[54:53])}; // @[RoundAnyRawFNToRecFN.scala 183:69:chipyard.TestHarness.RocketConfig.fir@237839.4]
  assign _GEN_9 = {{10{_T_188[2]}},_T_188}; // @[RoundAnyRawFNToRecFN.scala 183:40:chipyard.TestHarness.RocketConfig.fir@237840.4]
  assign _T_189 = $signed(io_in_sExp) + $signed(_GEN_9); // @[RoundAnyRawFNToRecFN.scala 183:40:chipyard.TestHarness.RocketConfig.fir@237840.4]
  assign common_expOut = _T_189[11:0]; // @[RoundAnyRawFNToRecFN.scala 185:37:chipyard.TestHarness.RocketConfig.fir@237841.4]
  assign common_fractOut = doShiftSigDown1 ? _T_186[52:1] : _T_186[51:0]; // @[RoundAnyRawFNToRecFN.scala 187:16:chipyard.TestHarness.RocketConfig.fir@237845.4]
  assign _T_194 = _T_189[13:10]; // @[RoundAnyRawFNToRecFN.scala 194:30:chipyard.TestHarness.RocketConfig.fir@237847.4]
  assign common_overflow = $signed(_T_194) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50:chipyard.TestHarness.RocketConfig.fir@237848.4]
  assign common_totalUnderflow = $signed(_T_189) < 14'sh3ce; // @[RoundAnyRawFNToRecFN.scala 198:31:chipyard.TestHarness.RocketConfig.fir@237850.4]
  assign _T_199 = doShiftSigDown1 ? io_in_sig[2] : io_in_sig[1]; // @[RoundAnyRawFNToRecFN.scala 201:16:chipyard.TestHarness.RocketConfig.fir@237854.4]
  assign _T_201 = doShiftSigDown1 & io_in_sig[2]; // @[RoundAnyRawFNToRecFN.scala 203:30:chipyard.TestHarness.RocketConfig.fir@237856.4]
  assign _T_203 = |io_in_sig[1:0]; // @[RoundAnyRawFNToRecFN.scala 203:70:chipyard.TestHarness.RocketConfig.fir@237858.4]
  assign _T_204 = _T_201 | _T_203; // @[RoundAnyRawFNToRecFN.scala 203:49:chipyard.TestHarness.RocketConfig.fir@237859.4]
  assign _T_206 = _T_165 & _T_199; // @[RoundAnyRawFNToRecFN.scala 205:67:chipyard.TestHarness.RocketConfig.fir@237861.4]
  assign _T_207 = roundMagUp & _T_204; // @[RoundAnyRawFNToRecFN.scala 207:29:chipyard.TestHarness.RocketConfig.fir@237862.4]
  assign _T_208 = _T_206 | _T_207; // @[RoundAnyRawFNToRecFN.scala 206:46:chipyard.TestHarness.RocketConfig.fir@237863.4]
  assign _T_211 = doShiftSigDown1 ? _T_186[54] : _T_186[53]; // @[RoundAnyRawFNToRecFN.scala 209:16:chipyard.TestHarness.RocketConfig.fir@237866.4]
  assign _T_212 = io_in_sExp[12:11]; // @[RoundAnyRawFNToRecFN.scala 218:48:chipyard.TestHarness.RocketConfig.fir@237867.4]
  assign _T_213 = $signed(_T_212) <= 2'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62:chipyard.TestHarness.RocketConfig.fir@237868.4]
  assign _T_214 = _T_164 & _T_213; // @[RoundAnyRawFNToRecFN.scala 218:32:chipyard.TestHarness.RocketConfig.fir@237869.4]
  assign _T_217 = doShiftSigDown1 ? _T_155[3] : _T_155[2]; // @[RoundAnyRawFNToRecFN.scala 219:30:chipyard.TestHarness.RocketConfig.fir@237872.4]
  assign _T_218 = _T_214 & _T_217; // @[RoundAnyRawFNToRecFN.scala 218:74:chipyard.TestHarness.RocketConfig.fir@237873.4]
  assign _T_222 = doShiftSigDown1 ? _T_155[4] : _T_155[3]; // @[RoundAnyRawFNToRecFN.scala 221:39:chipyard.TestHarness.RocketConfig.fir@237877.4]
  assign _T_223 = ~_T_222; // @[RoundAnyRawFNToRecFN.scala 221:34:chipyard.TestHarness.RocketConfig.fir@237878.4]
  assign _T_225 = _T_223 & _T_211; // @[RoundAnyRawFNToRecFN.scala 224:38:chipyard.TestHarness.RocketConfig.fir@237880.4]
  assign _T_226 = _T_225 & _T_161; // @[RoundAnyRawFNToRecFN.scala 225:45:chipyard.TestHarness.RocketConfig.fir@237881.4]
  assign _T_227 = _T_226 & _T_208; // @[RoundAnyRawFNToRecFN.scala 225:60:chipyard.TestHarness.RocketConfig.fir@237882.4]
  assign _T_228 = ~_T_227; // @[RoundAnyRawFNToRecFN.scala 220:27:chipyard.TestHarness.RocketConfig.fir@237883.4]
  assign _T_229 = _T_218 & _T_228; // @[RoundAnyRawFNToRecFN.scala 219:76:chipyard.TestHarness.RocketConfig.fir@237884.4]
  assign common_underflow = common_totalUnderflow | _T_229; // @[RoundAnyRawFNToRecFN.scala 215:40:chipyard.TestHarness.RocketConfig.fir@237885.4]
  assign common_inexact = common_totalUnderflow | _T_164; // @[RoundAnyRawFNToRecFN.scala 228:49:chipyard.TestHarness.RocketConfig.fir@237887.4]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34:chipyard.TestHarness.RocketConfig.fir@237889.4]
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 234:49:chipyard.TestHarness.RocketConfig.fir@237890.4]
  assign _T_232 = ~isNaNOut; // @[RoundAnyRawFNToRecFN.scala 235:22:chipyard.TestHarness.RocketConfig.fir@237891.4]
  assign _T_233 = ~notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 235:36:chipyard.TestHarness.RocketConfig.fir@237892.4]
  assign _T_234 = _T_232 & _T_233; // @[RoundAnyRawFNToRecFN.scala 235:33:chipyard.TestHarness.RocketConfig.fir@237893.4]
  assign _T_235 = ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:64:chipyard.TestHarness.RocketConfig.fir@237894.4]
  assign commonCase = _T_234 & _T_235; // @[RoundAnyRawFNToRecFN.scala 235:61:chipyard.TestHarness.RocketConfig.fir@237895.4]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32:chipyard.TestHarness.RocketConfig.fir@237896.4]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32:chipyard.TestHarness.RocketConfig.fir@237897.4]
  assign _T_236 = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43:chipyard.TestHarness.RocketConfig.fir@237898.4]
  assign inexact = overflow | _T_236; // @[RoundAnyRawFNToRecFN.scala 238:28:chipyard.TestHarness.RocketConfig.fir@237899.4]
  assign overflow_roundMagUp = _T_165 | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60:chipyard.TestHarness.RocketConfig.fir@237901.4]
  assign _T_238 = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20:chipyard.TestHarness.RocketConfig.fir@237902.4]
  assign _T_239 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60:chipyard.TestHarness.RocketConfig.fir@237903.4]
  assign pegMinNonzeroMagOut = _T_238 & _T_239; // @[RoundAnyRawFNToRecFN.scala 243:45:chipyard.TestHarness.RocketConfig.fir@237904.4]
  assign _T_240 = ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:42:chipyard.TestHarness.RocketConfig.fir@237905.4]
  assign pegMaxFiniteMagOut = overflow & _T_240; // @[RoundAnyRawFNToRecFN.scala 244:39:chipyard.TestHarness.RocketConfig.fir@237906.4]
  assign _T_241 = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45:chipyard.TestHarness.RocketConfig.fir@237907.4]
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | _T_241; // @[RoundAnyRawFNToRecFN.scala 246:32:chipyard.TestHarness.RocketConfig.fir@237908.4]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22:chipyard.TestHarness.RocketConfig.fir@237909.4]
  assign _T_242 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32:chipyard.TestHarness.RocketConfig.fir@237910.4]
  assign _T_243 = _T_242 ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18:chipyard.TestHarness.RocketConfig.fir@237911.4]
  assign _T_244 = ~_T_243; // @[RoundAnyRawFNToRecFN.scala 251:14:chipyard.TestHarness.RocketConfig.fir@237912.4]
  assign _T_245 = common_expOut & _T_244; // @[RoundAnyRawFNToRecFN.scala 250:24:chipyard.TestHarness.RocketConfig.fir@237913.4]
  assign _T_247 = pegMinNonzeroMagOut ? 12'hc31 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 255:18:chipyard.TestHarness.RocketConfig.fir@237915.4]
  assign _T_248 = ~_T_247; // @[RoundAnyRawFNToRecFN.scala 255:14:chipyard.TestHarness.RocketConfig.fir@237916.4]
  assign _T_249 = _T_245 & _T_248; // @[RoundAnyRawFNToRecFN.scala 254:17:chipyard.TestHarness.RocketConfig.fir@237917.4]
  assign _T_250 = pegMaxFiniteMagOut ? 12'h400 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 259:18:chipyard.TestHarness.RocketConfig.fir@237918.4]
  assign _T_251 = ~_T_250; // @[RoundAnyRawFNToRecFN.scala 259:14:chipyard.TestHarness.RocketConfig.fir@237919.4]
  assign _T_252 = _T_249 & _T_251; // @[RoundAnyRawFNToRecFN.scala 258:17:chipyard.TestHarness.RocketConfig.fir@237920.4]
  assign _T_253 = notNaN_isInfOut ? 12'h200 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 263:18:chipyard.TestHarness.RocketConfig.fir@237921.4]
  assign _T_254 = ~_T_253; // @[RoundAnyRawFNToRecFN.scala 263:14:chipyard.TestHarness.RocketConfig.fir@237922.4]
  assign _T_255 = _T_252 & _T_254; // @[RoundAnyRawFNToRecFN.scala 262:17:chipyard.TestHarness.RocketConfig.fir@237923.4]
  assign _T_256 = pegMinNonzeroMagOut ? 12'h3ce : 12'h0; // @[RoundAnyRawFNToRecFN.scala 267:16:chipyard.TestHarness.RocketConfig.fir@237924.4]
  assign _T_257 = _T_255 | _T_256; // @[RoundAnyRawFNToRecFN.scala 266:18:chipyard.TestHarness.RocketConfig.fir@237925.4]
  assign _T_258 = pegMaxFiniteMagOut ? 12'hbff : 12'h0; // @[RoundAnyRawFNToRecFN.scala 271:16:chipyard.TestHarness.RocketConfig.fir@237926.4]
  assign _T_259 = _T_257 | _T_258; // @[RoundAnyRawFNToRecFN.scala 270:15:chipyard.TestHarness.RocketConfig.fir@237927.4]
  assign _T_260 = notNaN_isInfOut ? 12'hc00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 275:16:chipyard.TestHarness.RocketConfig.fir@237928.4]
  assign _T_261 = _T_259 | _T_260; // @[RoundAnyRawFNToRecFN.scala 274:15:chipyard.TestHarness.RocketConfig.fir@237929.4]
  assign _T_262 = isNaNOut ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 276:16:chipyard.TestHarness.RocketConfig.fir@237930.4]
  assign expOut = _T_261 | _T_262; // @[RoundAnyRawFNToRecFN.scala 275:77:chipyard.TestHarness.RocketConfig.fir@237931.4]
  assign _T_263 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22:chipyard.TestHarness.RocketConfig.fir@237932.4]
  assign _T_264 = _T_263 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38:chipyard.TestHarness.RocketConfig.fir@237933.4]
  assign _T_265 = isNaNOut ? 52'h8000000000000 : 52'h0; // @[RoundAnyRawFNToRecFN.scala 279:16:chipyard.TestHarness.RocketConfig.fir@237934.4]
  assign _T_266 = _T_264 ? _T_265 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12:chipyard.TestHarness.RocketConfig.fir@237935.4]
  assign _T_268 = pegMaxFiniteMagOut ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12:chipyard.TestHarness.RocketConfig.fir@237937.4]
  assign fractOut = _T_266 | _T_268; // @[RoundAnyRawFNToRecFN.scala 281:11:chipyard.TestHarness.RocketConfig.fir@237938.4]
  assign _T_269 = {signOut,expOut}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237939.4]
  assign _T_271 = {underflow,inexact}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237942.4]
  assign _T_273 = {io_invalidExc,io_infiniteExc,overflow}; // @[Cat.scala 29:58:chipyard.TestHarness.RocketConfig.fir@237944.4]
  assign io_out = {_T_269,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12:chipyard.TestHarness.RocketConfig.fir@237941.4]
  assign io_exceptionFlags = {_T_273,_T_271}; // @[RoundAnyRawFNToRecFN.scala 285:23:chipyard.TestHarness.RocketConfig.fir@237946.4]
endmodule
